-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
f9Ot3le3rJihxtkkXy+5BUDEPfciT8HUArMHtz8jRadGM6tC1S5cf+Hbxv4Uqm9r
1gsqubXsyfL+Q0xoLU07/w7Hru3+tuZOuO0Gg6mx0m8yu4nFOlTh24B0M7CaPNmi
OX8cmPyvRNxZZ67emfwQgSRu4BA2ScGf6mJPae4zC/o=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 6496)
`protect data_block
Pm3NZKKSo/Xl/vyvoo4D52q9fkB1spgvh3IW1wocrCkcfeRVtl1r8SWZDQ70C3i4
irjFyT93z3EhulanendfCeH57wobDKgnX+UvlKKBVrGAVvS1qsCRmql7zA3FynOS
tXRAdpYUNkZOVtYa9FAopoZjWzfIeYYESeglZA51khjItkJviXomHJbn+Ls1VBVn
EIiKwpoMD3BhnneToAXHHovm5kgEY/SEv33X5qEVGTE+gNNMn90CX20K/oGka0pl
PLg/8TkAJIuBfnXmzG10k+KL+D5InNsTd71Oz9P/qOtusnoOfXTXdXw6SE6SHoXj
0riA/EfkBmQWt1SkXL6GaGsSI3vXz4y94DFw2BErDjh+r7zQrPFFUgdzESswFD/G
sVHLxpG6pJ53qllZLaBl9ChJzyavArWEuV1M8XEY75S2GHOqeHo1BvkIzZxWxy9n
UBcLwM4bRXN01Gb/1L3QgSYfrVu/HMbjPEHuS2p5MFjymhw3mgFpYXM8JlZ70Uwq
YmsWpdvjoq3i+UOAQdN26R9ytslyoxjfuV+DZ2pPrNR8A9B2/HqtceTKiLUvpc+8
dzMNs3VR2TD6vvtNFtqQVYrrxY4iVWYoBy1esItb3+zRMVDOcO23wv+By4e6hcGw
2EFEJj3ul9vcUWUVUddx3Is04bTXk4KsXVNcCqz8fx4yrQXrSGMiW4IYwSp1P1sB
HlOLVnghAF6rT/z/fGyR3XeaRPC8061j/dpg9BYpuZQv676WCp7ElHgFsDF0u41b
5bj2NvQuQFlITnRFw/qOriRyRNOogrX/Q7bjevbPN8T2Istlo2DAc363q6eJV7Cr
lCXPNkkvFJnUCZN65C08gnXIiow9pAGPhWWURedDvaOWFqTTgETVc919V6hhCbcc
6e37KLo9g7uxmdEPjPtjJLpx9431XZLh0ssfKbCEAUX2SPggXt8MoaCDWBR7SFA5
ducRWWwo0TDw0uRb0gWJVtP8IdDLf0FuwOI3C+PEilKw4VXO3USPtTWquPcY0yy3
k/l1pVVwdIPtYjWgDSKcrxoynEDJ1SpZHWztt5KudDiiJ0q6tXeKF2MiTFreDCZD
S6AYuB4XZ8qk5mMrJPoCVYY0GB/qc+xY7m055Kl10F+IdpoqSPmyZxHtGcxCfrxK
Y9k3YbYB9zQAcJiHunz1wV0Ew4aXUpwr8/hyHqimJ68I22pCgXkvyKuEbkuR9Nlj
EXjnVZSnlq7z0PtKkamRMhtEt3zhqMuI3hXs0loqWt2Zr0tZI9pCxHbNcvpqA2fR
0mfyycrOm2Fp28GY+0ZqWhcqB9ozDclHrpJ+lk/rWAN1TIl6DCGx15CwGDWfzxgc
cZL8Rp6f8oh4dOENDFzTo7aLMjHAlBae8WfveQ8YzYYBIdDOLBe/gYA6C+HHV3nP
xb8qq0fWle9yRUpJutloE8P5uE7uKULENDPIOBDMaci9ZlzUFTjo9UjqD0mE+L6U
bhYjM+41baJG/CGbuUaLcpNVfHU3Z3d/8PW4go7zT2Y/63ucb8wuMfXzaF1T19Vj
kv5UsN3OesrL9y6bt8VAYAjWYPoB6TpMeCJGyIoQq2pzHcpFGYkTray6RoBVAYig
+LfJTQTqyRSqBDjkLC3dYY1DvMhydv4ugjPGmQc/u9yOu1VMDV3AWfDgIR6B/KOT
drTzrF/yuNvbFlmOkNrpNNdmYFkSs7Vc9kyuk5Ssg/HRo2J+bgIaS45Tz2Za3BbF
VSoa3giqmTl4j/miwgjTKLrVp7QCFm31thPUJUAIOHcyIvLFeharzuke0UycHAnQ
cLF70Oo6ht/lMZlhm9C1FRUSmuC0m8TRQzTieFl79Jop89vCdlEULgvVmQe80BA4
yvuk0wIm9J7oomE0886ekqlt5hzWAQlj//a/QNhhjvps+Us2QJ4HnJM3I5wjx5hl
9JGj8WPCwxpnsE3f96Y6QFZgY4Lw3xBntuuzIZofvcL+5Qbg6uh5ZWNqqq29cVyp
7oFkzfgMx4OcnbcMu2evQYZz82QRoBHIKAl8AB/KvHop11UuVx7I10EpeRK9BVJf
lyu3yT2yMg3QR6+2iJxI8RF1bud5uaxX1PMUmmpqVIF4d0JwxODob5lldMdOdys9
tqo9IqZD/s/brIEKQu1dwhI/AjN7mUFlD+I6l/LZnGhRi5WRuRWnO3mb0NhNme4O
28CBkYyY0W3W174YPzw7vEMkZ4bxXZW4nGVTh2Qk4A5pgZLN0MoTXcb+kHAX398n
QWRYh8JqLLL5ZAEmvePs+JNKunv5Nn80d9O9GewJbBzaMhKpM9H+5pBmQ4lHI1XV
n7kk6MhieY/vEVnr4J67JG8pr8xIm9RFzGJCxmyoVWoPVbLAXauNzO6L5oXBGbOT
AqYdBZG/XCKiMTAPBHPLzoL9+XGJIFDRC3GGdKak2lwKGBVrUlBQaN6i1Bq70+/H
T7bdMZU9dtEMTYDKdyUfONgka377pvG3RmXQ4DdTZhzzkHazRQ25vj/O+ArAgtKA
QD8I3YCLjuZRrjwG4/9/GwLDCzY3WQc+B00s7lXCum0X945+W/JtmZ/2DuUSp4Z3
aBKvoZOft3POcOgPqdeHgcJ9qWrowevZQ0YLZzPloqRnSvbguPdz7iP7W7WbpD6c
ksKOJa8l6qZFinxv7Vxfk441BDGTRedhStLHJA4Au8N1atQsL8uIhcOK5ps20J8J
npZTd9spJP4FF11fgJrtolAKe53rUZoTuQJtQF3NHN1r6MIFEpcOjtwe+bxz+Oca
FvmlFC5yP0toRpF7f9faN+RR6FP0fxfFs1Otjigp04tlxhGzWSQq0UI/JOE2eIds
usQcqdY31G915f5lnz7mvGoG65j0mWhV7inzYzXRqrn/R+KtzAVP/yjaKxWs2U8e
psmrJIlm7rYwiZfP5G1kN3TayZIUzG0tadXHHz3zgVNTMHVWwtkpAGeoY9JTpr3G
qlGyU9ZBsvZRGDYZ5I5Nggru9VILy3C0VdfU40VzmA2cBd1yWgmVHWOlVMvJvrbx
GxcQEYrg3gn+tP5ceQuPuSaZ+JKpLhftS7tIVyJ7WNoi5XDxj/Se+6C0eBxpyjUd
dNV2yU7Vz5Dr4Jyppu+oVZU0aenWSCKGOuIyDV02nffzeReqI3oU1WOaAbQbloyV
Pt9Ta0P0vTZgklp7Jd7NyQuOUh/jOULKEn8SAi18Bicefzsk+9392TZTkAmd5SpY
DBqo5n+JI4ks8w/5hsb1slk7rIsHfHpk/Tg+H0bdgVWpW6D8nSGNQZNFlXW0fr5C
F1y9+Atlp/6iLUCHK9sTj2UcZlR/0ImIvom2IoL/+3ZR6W9mxrmZ0IGdWlhgzcvj
emn9PxEuazdmEJVv9wCHtLFWzQLpMwP+niL+HDbVQZLiBORT6FB3c9RYP2GCrRjB
HC9iKiWK0EnQnfcmU8FaGg7UP8n90Kxp9GVVvf2fa9j+bHMHvKW4GWwe+y1AWy4z
8jHLBkluSr2WMMQR6sxDzgrbckd0uchhdlzjItC2oeD1SI9/dm40qujLRDk/QVxZ
nMfD2jMnlm7ddegq+g+eXy1ToFTX5XfqLsZLKaB9Hqe/6cBdlTIWyrh1oT2HBTmi
GixTzHOXa/HCpAUFZ8yXnPiIh9XGgLz5bmmjf53zQkn1JU5bUFQEz1MzyoFXLlsf
axZdEivOMMuFynN7J41t66HFjfiyaR8U12F2461qNb4VriqV/H+ks5ixCf69JAQY
g/dqB5Iw231W8UXwCSgSlOGUM0hc5gfVhsjqVVEisEOShfuFnrzdWJpaCL8N4C2M
7S3syvfFAtr3UClWLXzGu/23bvhfhgb2AoXS4ggsFYCEeSZhkGy5S3h1CCNMBGl3
dzYVyqJWviM8qpx7NxfNeXaEiiMAcpYddE5EIazCMlht7SghSA8j94puZCrx7Ma9
yFglIGrNhDuszvvqPJKbaT+UPCO+dBTo3rSNodZorfmCo8IO4GG5sRIq2fG96FjV
TJU/CZ5sAn9N5Iol2lCvv0I9wFHns24UcJ73m+yO40cTHj+cqt9wK1XXgs/vk154
xeHUWPzqD+aVtVFCfem4MtoLzwEOFWQq34Zy/a0dWR7KK4l5nMJN0Xgz/5Jw7MN2
Ei1nW/SoOWxzRNbnnwjBDeF3JRN2zLs5MKDbmOHPFeO+dR+ku7reSeeJvh519Fm5
8yyzDoCFQd7W9A9IMKoZXc6Xz4kJqf8kZUC7DLUjpF/b6csNs/GQ3dMEgwUiy0xq
arSY+QJAcMMFkeTE8by8j4yM4Amh05P5cva0869iZdBzLeLgSk8bs8BQXTymi6zd
BFp7olD/ppCsczzH1Tb7n/BeTbK/MhejxRw4oGNBB/SLuJALtnIXt7V4efSQVZLP
Ihc+FD77ujUxaeyoOahccV/wXo8e9Y8a1N40i6BS58Af7IEQ1to+fZn0eCV4jWS2
qsKSYRWzQwZxtuyvQZst8vcCGQ0UociNP/FH5vlGUqT4+qwnBUPsKBIjwQmI7VeM
g8kKLcCMehf9e8xAvfD0jL+iUl209fWNaCzcenQx/NnieZZgH/nZZ1P7O9hyOnvV
y2Fb2QXfe7NOX3VJlyxTJfykk4ld6bpYOymYU2vgcz2VHfXP6S23545UCJy3q8tP
H1t9dEHEOLJbeuBkKSqGWlwjr7emC7DebRkyg13PPJBno4iZM/vUt7O1nG7F5gn3
9juORuTtjooc34O85jrIVVDlCx21PouUK1vkNaeh5JKiE5ZuniMrnqYdDDsSno67
3cQCa9kpeIhdsbWWHkVU4ulyzAxKG/wUIHRTwg+mXq/2rMyvFUo/PE6tUq8HTUtY
FtgJ93BzCsB3GoSggxDvJZXnhyn+0L8qxnAFNvGIfoVpbmI9p6irSxHXE+MRxnDm
lkJdI+OB+P2GlFjLoWktcOSuxjtonbjkpoumKYkx92YtII30An7O035h/JnHS0of
PyRCDc4NbFeQmjZynOM2wZvO8rWZ9nwGyjHxcBUbujqHSnAwH0NpuYR7pJiN21KP
Ltmx8xD/eqy8/hNeWwWFpwYjAe+PIRAwtnmhBDeTJVGNcAvMdIhDdZITr9+iXGhz
LseyokDEeOVzS6WTFdLN7jyg5NuKIp/x9hL+Ssk9EDaJFpZ4jQQ+SxH7CEVGdTNh
7TP4JrVkmGaJMFaAcZSt6Naur6gMg0IAmDVRoPbUwIvD/NjP/0ajmMMhErxSESqx
vEYtMiRHuG++wWkv2aVEWK0oDSKUU3giRGM/x3kN1ds9R/KF1guD6+NVIHVWUOPa
lD6K5YRiE69AJlANpvhBVNZWgIqHYuTupOyN97sWBv7YSVfRVJu5572ojNxv7RpZ
bs5yOuAzm9MMhgslVKEALc/qrwtGY+WQ6CmG6vJszN9tOf7hIdeXkFxsP+9zWac6
mn4opvKxwjPJrPavhtnvNk1W557y2DcKhAoP932hvFBcyhRhHHQ0s/iIaNhmzD15
Rkmni3kh9hCsGPMmwbm2NPgguC5fg8u7RFHU6uBqLvROXwK+sb1bFe2ctV1nPfqB
DTC0MS5aUh65Yh5sO+SuY8/VUHBTnRA/vxn5WtO6lZBS4Kkc8t1gaHE29xRK1j1R
5dYXOehLudzHSdB7Fo1SyfC2lgpKOtBUCCrNmCGRtj5T5BXzYALVfdC/u5LKMGio
0S/bVnSEGgW7ytO6G66R/MC7iCapfvR0poo3AO64iAccRwRBCyeeVkeV8Skebh2b
3o7paznnGMwgixNI9LYh3ghs6irhJCDFsBYn1Z22jsST1L4jscOzb/VOACFTsp09
7ZADy0WOT7n2TjU8MhqABI2FM2LtCNAG1oxytrgNKMq3nvx/c4zk+NGeS2TYJzzg
P1cetzHZOnr/p1WWyJLdcZrwdr0SY1TNmZ+/kZn+DL5OZbqb64G18aS6fZjbNiPg
0nf0Qxf9WgbVdDHHYophwvyP67KJ7fCoMrYfOJRx9s8BfmKnq5bXslG53UPFheOU
pNJsOZGDEWLBBjKpgkgxMls6J6vQhTUzzk4jy7hPAyZ+geHcqpfTOF5mTKOIeom1
2JT983zjSAnAcWXembVTYZFPbLYpWpAIwLz0rnFHXxj0Zb5WpmQm0TYyajSyRAq2
CvFrhepFU9xYMVCUnUg9NoRbc34E2urJpUfLTHD4kSk1m/wIAKjm2oTu6EzeWi+A
Mk1+0ooePeU8qRMprDUMteF4GqXdUiT5gwOCZymZhf1hHHF2JfIViYvHgSP0Pofr
lfsiAq5oXlq2Jwle7TkGj57s34w2WCA8zr2G1UUO5U18wELdyRvi5PM5O/Fp6NLT
CGvtTUSbsVXOH3HVWryRoNiJLkxHLz7xLoQ5Ki7y7oI21WZf8hR8PgSx6+gE0OT+
9E3hqQYetqANbHmdCbxK8mZKn6bx7aN2q9QO92/wwqMOkDk508WrLRTwFF5phMMk
xO1yOgiIRldznAWZx5MbO4D2mpVfruy7zFvbjZ/lSvkp8GcJFf9BoFHKF3kYM0Fq
G3bepjNa/4X+eILhMfnQmJek5ZUWvNsfm9kiC68rHMoREY8gCoby5E5TzPbJsgke
4ZIbpPVVd+6N2CbUz3RJ93vSv+MQnRkNgwn5fyV3vuhorqVpcmyBN3TvDLLRqmtE
huCVJxpmZi1aU9/oC3toHM3XytqAyB2yM1eRf9KKPQ8YLVRYOMgHvx01B/hvPRjZ
Cv3H8g0NcC7wRL790+ephJ9+xYbn9LGtisTrYMIf4rJQ8zK6NxlFGoXaPlT9x/ES
o+JA8W7BoPm7Na3V+DpAxSjYDT162r5JISUia9ieLDEYqFkla8kxwWUFO4fD8DdD
OPgEOZ0Ad2dytnPQ0a7uBTDC/qTcHXgfx4jthcn9JiSI3YbdaMVm/5NeMFEF+pUE
r++KYdD7PgrtCgYVkJeBZWSMBFS9qc27GPyT7nQf1L9HSwsGGsZ77hBxiJ/u9M2F
oWgHeE9sDsDL1zCcjR/1GZVb40cotgQ6oHxAv60BHfo6NqeO7zbKMxy+ViU/rwYj
K7Nfr83JRSnqxaN0P8inIUQwHCj3V7g+tc+sLaIW+tzvWj/MRTX5P1alwcaoLdgA
doTKA34ZoT7TGiG6Q98fUxcB0gbwv6b1okJ+/XViPm15p6YVW8HSxE8zj9qEsxoU
VQCeXmYMiEJpHtEY+oJXLxtAm1cia+oIEiIdaBNZT6piL5IxaTfFFggLLLhI8eWj
wxBqUeDfTg3qHPtis1YBntNxa3g/Oi5VAyrBX6E4nDo6qXKIzs512kcaff9/Pwkt
PrifNdkBhxC2aA83wV96UqGIgF6Z7IK0TMMDtHERJ5W7ad74hqCbE2cgf7RjvSvi
9JvT6DZft2EwBzcVAv24+PKVI1O5fOh7b46W68Pk1zI0PTU6HODXGIyTNEVRMqN0
Tk5kIys1wQbczXbXfcm1/d09bo8sKEiKM4+i7CsuJ1cu3ZYrQrGwtJtb7wWEdkvR
g/+C0SEJdg6Qo07ZJvTGeQecGZmhWFiH7RzN+WkBdGFIUaupYX0BSO7rFTRuLzH5
uV9HCzcrUK85AJrTvkcknMcsIBlnLBOCfSEAAF0B9w+JvHG8xaAFf6JtFVuP1ICM
+Eyn/tnFesmC/u47gydMDsFGDwcHb8dpUl24MjGUWQHS6GspMpppcUHKrDIxMoLJ
/JY60PJzNzNzPtOssTtY+54jSA30PLPAIE3PtoXZjJGSKPo/iRPBZ53atHYiKfgk
wWtgxxjLA6CZl7U630sURhB++xCCCzvG7iJ7ouwvpGgTcgxmsspjzmqpaU4tWZq5
qFha8AU1TFDDUIRjuSmrmL/OfPSjnWUbtsJxEPxO3TCfSOjgSXxBAi0QTFA035UT
GvNh9dRnur2rb8wLabv0Swo262rlfYiarV3A78MMiz5/0BfV7Ea6HBsP1a6eLa5L
15QazDzRbpXyYynrQjbx/ydx1eO+vAF0ySb7RORblhw+0HEaiN4UVnVYdKeRklih
W/SG0recwQL8cZyMIIwfWZWIKp+rPBrAX+pw+Go9cx5WHYbt5tKNsFX6ntCcX5Rt
KhnrFK7qbLnUs3ie2IkmQRi/7uyl00IJ0IkqkgcNtj9NvaFp8dbglcn+f0yAnn2i
Po0swtltBtd3PN2nHp20AkpwfBh6tBg1jf/za6GxJ3rhpiRMHkFnOSfpwG3McZT1
Q5g1B3mZnbnnEpnsSr3hwu+MMDCO8NUPfp669GAwebc9EuqxCnPg6FwQWQ6CXVXH
lRBpBPhqGeapZaWs6UneLJQDH8SCE9uVFY2YUa8g/Cfn2u8jNRbXzpwoPMBKFDHv
8lnAkGjik6Ox12QIYl+cpjbAyuWJQxvxA/TL0yvrRGfrgTKpLJeSb48z7wtNUNus
b3txHjaYtbLpqhZaMZ4+Oxaa5vWQDIsFpQM7oHOPxwB3my81Lkg25/41MuMRoEz5
dHsMeoh1FxWSH4k0yJBudlPob5gVM8fQoAGFgj3Qu2CSmV+a3Diw4d6ZNfr8MLAs
SkL8pEHCzdaiH7xy1Sc0sTZyooCvb+n6EEKe2ITkgaTO8FQkSCnpArcaKsidUSDj
YO18uaqBCtSczyzKRibGCXaSPMfc1ILSrEaHTCTb1V2tu1BxOszDeb9AFSAikHqC
9RlFlJHOuoR9rZV02hIvjNnHEiFuodwA88HY0drPSZ+XX88JTPl2MQsSbrKHGkpj
1aHW2nggfD93Ap1Qx5yiWw==
`protect end_protected
