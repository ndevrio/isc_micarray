// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
HM4@NTWV3<[ ,:U TE\:5GEUHH>!-E^']85ZN/;].%/_UF+/O 1W ^0  
HO:;#"&)C6SRM^VKUK;9OI>)(P]1-=0;#,6)2-&/R]N>-1P&UI0'@DP  
HRGN,)5;^.>_BM%77KCQU)]F)-@X0N;:X;Q+0ZZ4=AZWFL.B48 %8P0  
HJ0 RV+86.O?'KB!&]4F(P:Z^#%OY\:^?'E>CUZ?DOM-MLKQR? B5Y   
H#B5HO-U*"<3)Q:(9W\N<)@P"5=CPQ;F=A;[!R9_+HRPGMX'9,@04>@  
`pragma protect encoding=(enctype="uuencode",bytes=13920       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@%S0H2#&T=F53JG-?.-_WL/T=]&;2RZXB!1O-G&F[JUT 
@;!S<^'D-B&(+.(;;^TPJY-^(CLYQH5^U<LGJ?Q,;*!@ 
@XS<0$KBO>FP'BQ@8?'X=\ +=T2SYJ4 N7:CB$KU;KQ, 
@.5AS8IM@F/H19SE1B%,D<('*'_,$R'<'TH.^?8#U=C( 
@+R9>:EQZ]PPMXF=68N.UZ9%[W][-K_CX&#G$+/VH;I, 
@>R-8:*<8@<C(]!!8!]Q&!:895F9Q?3/ZD(^CV:S1,YT 
@U(C%:A:YTHI$V"8(BCC0]+3^@4N:!$#]7+'B'-!"95D 
@P! Q'V*7^-Z,OD[YQT)/D<Q[A2@EZR!A 5C+$S5 '%P 
@>G1E()4::YXRO"#)%I\52I\N'X'I=PK'BLY!>6:G[5$ 
@M(&_-/1>Y2JG:.]&C8[>Y=@2H^C7O+"+7M+"Y-X"'IT 
@UX+_>1PF^WV1=US<CBIZOD#T.B O:3@:K_,?KU<'I08 
@RA77&::=MW_<N#]Q^7-4W/X*JUKJ>;*C>%_"MF7"&*\ 
@$?1P"A-/9D8RG!*'1[.>>AA?;537/\B)(YV<8XS%!Q4 
@Z[VH0:NN4S)2O6"6$GOXM5FIC^09Y 6U[\5],?]UWN  
@&Z.EW06;FZ_W!HZNE+Y]U A/$V9]K[YN/S;!&!:G&Q, 
@<]?FDZ0!O\0[7SS)K]M2[6_\F#8'&,+812-JX$$TK., 
@T<- )1Q;D/L2T &(A^:U<Y*H,\0IT;"H$F% .].BA7, 
@1%1-2O,&250P&#<CXP:G"Q>CJ4/L?CK=B7_4J5K<O1D 
@DLA5+QGF9?1FGB]8[8\>6=%G<QZICZ@A<X%MB_//CW8 
@-Q'WRM8WCSWI6MJGLIZM,3<\:O."/?%MCDCWU:1;DPX 
@W,4F.,S]JSKA)V$<>2"GYS<!^81^6<U5+-\5FA@N6IX 
@:W]BBJD4*H%&4R +#H4FYLSN"L:5HM<4L20P[:TW]W( 
@13*1P/)46AC*<,$2_^$)WWAG%_O#[=TW=\4&VN9C<^( 
@0I8Y[BA(,T#286)S+@/D7!/:@K XT<:)ID*+R*E>(E, 
@S;5$&8*)I-7KJM9HAB)4[P<]Y6&?I%1J$\5:\I\.G4\ 
@=T*A*K/$K",7=A=43!'Q(8(K#&P_U5+/2P$O9$WJC[D 
@H#+Y6Q_Q6M%M&JA_=G*'1K3$F#57% YB D9B +=0L^@ 
@O#.U"*_Y,52OLUJN8B-T?H#GV,\9I0 F<T.O6T?::7D 
@W8AGH!JY7V*K= KQ$9 II"%.\10JM9DHEY2S:6\"AL( 
@\5'7-+;;,HZV-&O&(G(IQ0!)X]()R^GC4YF_EWP14.8 
@GESP*D)<T?4Y@>VMX3M:@! :+_%Q0K.]  CUC84*5"  
@<"/10M^#?H!"T8+I.KF:H51*$:95OQ8_A< .'?COZ8@ 
@/,E165M)H3^$T<F7?[MV[JQL;\$$@QJ =C1YNAJ([DL 
@"S_:^PG':&Y?Y?Y$04L%GHF+?8D18EH@5%4$LKW@<QL 
@7R^1,U,^'+;!0L33_!7PE<G(KR&EH!%*=-]X_]=1RQH 
@7CGC%#B'HR78] #W<I?NPF*BL_=O2CX)#%2":KERA 4 
@3BT'4"2\3I+"N0I->_CDY!8+_4B*Q^H7& 4RGZS6>V@ 
@*,MH^[-/W<<@7.FOM%I%F>:'2,\L"<!I)2=SNF[@,18 
@!US][XI!<5J?GMX)Q(F!HZM^-PY^OO4O^WRI;L\*8A  
@/KA<W">5).GI N>K64NJ\!PPA*TE7S"?]I?'8"S>D2P 
@()JWKPDXFF;&]93K9M1<%LM."Y)16(ZMJIS6X\P[]%, 
@FR"H(@OACR?PH,@H$%@XNW]+DV,\^RZ4M[9YV'%-'"4 
@@)9&P.I\,54VV44B?7E=^ZHL$6XM:=6>YJ#8E,20ALH 
@?P8/A:/</9\N \W3.D]"DDPX-[3-P3"BU(K9V"2:%?D 
@:6]HHWXR8GOVA>K<'0J@'*$^4?+OVW3DIZB.$>@VUMX 
@LQXM[T+%5-MS62TLLB8$'<8D6E;<2L6=6UOREF _R"8 
@#-^M9QP@G;F@[CSZWMN\/#?0F*1*C.GU0;"TQ0:,,*$ 
@NHC2X/6$P8AAE=:)//0\'9^) Z2J>L$E;N&:+Y@MB[, 
@EAXJ!.%_ORH>&-(&WOD::7!N&S=*4N4DO^W&3[1>8R@ 
@'=Y'G6T+ZS=S7B\N+4 [>K;GVNC(=CK-C+@DXZM85-X 
@$B@1[?FZ2M_ZOA.'DF=G+XSG*H$.@R^\M; \BPV'HGD 
@8?Z^VM"XQ#$/<=<XP)5UM4'_EHMJ#27,^$,V&GQ57G$ 
@TVALZOTM? 9=$HUQKA"LX\K3.LI]9.E VC.-XIN$,6T 
@U[557KL0D5V:^T(=G+X3+P4G&VN]Z+4C62[XX1+I^ZX 
@A&@:96XD/IH0<:!)UK2.%KMWMZ:3U3M>L/C-D,!8+60 
@)JO+8R-!UH;^#[0%]:J0%L+*O:MDKOF7382@CSG,_'T 
@D1GG3F S#<D8W;@<MK*6C?.#&YOW[8$3&X$4AN2G"H$ 
@VXCBJY-S%>/'1Y^TW&%323G:EEN(X:SB]RW.PLI45!\ 
@D3$3M1!X#E/4<WT>+ZY;@D_7H'P(E9*\@ZCB'=144Y8 
@%1GKEYZ174>6*6[? S.W(Z[,BW%:OVH#*W+W 7ZROD$ 
@IM,E=X R2TDP&1%&HYI.4^,[&'\\3Z4GUD,>=5XW4KL 
@]9B]H(1MHRH9S^H(?NJYP ZN214V6VX- @6<E/-6:', 
@S'0$W=^26>Z5<%-]1T\W<B1)T0/&&SX-[+]-!AYC9R0 
@C'$^&#^IM GFMW*(M1!0SDB[Y)WV= QT7(\0I9ELJ6\ 
@Z.:Q))2-&U*RP]LCP]E-/7ZZ@_"G3!1,YH_?IO;0G,X 
@4''U!Y+FZIEL,F+C;3H]*P2\%^R# $8U-VQ"/3R*C=@ 
@M%V:75)#CDI!Y\T8>;1T)H,9'/4>WHL^73HF(7=_^F( 
@SS;I#F8;+/E(_@[/94>J=HOZJ<ET0:\-AQV*(.VH&-H 
@E .+>ZP$/H+USS[\+TPRA^V'3R]]3=J!*6;2><YF&N$ 
@I(@@%;A25^L]"LJ.J!9\I.#QR4*]EKD]3!55VA)=OK( 
@,M>X,;O8+".Q5/,QW59E,F^?M_&]NDJ/G:6?MBS(&G@ 
@X5F*O^!D'&!3??JQQG4QV'6#C1YUY92%\,F 8SI!]9$ 
@T&W9?^U*$A[C:KWI2N,R/A&I78#WS*]W)1I'.\?&C1H 
@Q;5@F@;^"TK45.JB_4OGHTM)"%O[M<A\I,\YSC2B 3T 
@\3O7WD)#2A'[YO3A+DF@@C%4CYULW7Z.%;H\<)/RR&0 
@'U L=G/=T3$16]/.5(4=,*D)1I?4L!1#@5L8J)?/ZC4 
@!11Q,C[/3V^HZ<+;[JHR%]6U/VG7R/QH 7I>9Q 4?[H 
@PG\Y;;@ %V?)+.W?YCL_!+Q0H:(!!&P_(!$L./&43]8 
@%(. )N\@QGDX'@E OK\%.^(<8*8C/7)\^K?(%;NK&QH 
@<&"3;@J']-G'MSO/<E@&%_4G_&B/L09&$0;GFKG#Y:4 
@];1P@Z)+\@=L;%//.4X%,6)4"UQ 2BXPU)WYQ67*C[P 
@0$/O.<>>W_'$ RP2U+%,&AB<]U#H+R\C/$IRL<:0FRL 
@;OAV6Y#B,WQ*DW]\O&'B$MUROZ<-@"T4CM.W!G?4&5\ 
@35^+I)T12+!&?J^4-*;2Q^L]!.?X)MG+1WG3OGA+M*H 
@K;HOR7$V&ET"I7TW6K'$TGPU;=!'-$BB*5<S\_<1 (P 
@NV8V&.9K-W:'LMO9_@@\#UQUKL(7WB<+OO.9V#-_,,D 
@-=J#Q0A](+2P7G!A*)FR0%;G^*?:P")4>O$6^1@=B9@ 
@L0N\S(8VBJ2_B)IN?[LR0&B'(L">_=@MT^^Y3J$<6SH 
@8@$MU1PS<&0H2)THFS+J[M%:9&$JWN3VXOI *>8 @7X 
@X0DCN3L%7I:;RM^3D=28S7L\DI=6H( F 3'!WSD2V9( 
@*6D1/BG M2#4VEUK3E);_YLI&&8L3KBL&X;(K*_>L<4 
@21-4F<Z+:D9ZS[9S4N-;AU+&S Z_08Z0^60EWFON3H0 
@Q[]O1J@.<-)6UCOKG5F][&J\X7(6W\)UETY-+N26^X< 
@(4<7>7T9ED  $I:45I5B@?#$Y* $X%-\^K9IK5.D0E  
@;$]FB@N@15Z_,$([STIL[!%NI^7V.0( ACQ:O=C@?'X 
@''SCE=WN$3!.,J1A\ST_%UGM/^])9E]1?H$'-)RS=3$ 
@[7@+(*?XWL#+G)\ $@0=<D_V;NE<M?_\DF(JAZG5SY( 
@&+"S''ZD (2RZ9?_L;A67R[?&XBJ#?J_4IMRQLT]&KP 
@,'\2?K MH%J-5^U2'/,@@IN@4G!%Z+%^+%!@FMS,<_H 
@X%E'CR&N&L&M!A-R%#GZ!.%P2OJEPSWVPH1[2G/1NP\ 
@>LP4 0;$W"0W9M)D:!A5*&:,>"$MUNHN/VGYE*B7QZD 
@QP[!D:PT=W%!VRA*'27?Y=K9DIH5$6;4X709A9OJVZ$ 
@<! UR;ZR@;?*T@ ]$K2 ^NWS6=@+-R8/9V-3=/-M].H 
@"H]51NQ;"?^(C%>OG TLVJX#,LHC)[#&0JLPFX<I7L0 
@V!@(;SEB0 JVQP=$.K@C?Z&$G8(YN -;)*JO>^3 ]YX 
@,E<UC"P'C.#M4)Z2-4"4Z0:.?RZ;UE=<F9*MJ?H_E!X 
@%O=QZ_Q*;W]X4QAAD!A5OT+)('\P3"V(<4*:M(D&7F8 
@6M!*_=- 27W/<(#*2! RL[H&-';F%_Y:EMEB7ZXAIF\ 
@PZW_W3*E%O<  4!"8$15IF99PK4D:E^C+NO13LPGHI$ 
@M*QL]#R (5#N2(S/B^[?=ZT&BS4I2%CMO8R?6\LW==P 
@..Z"[E2-&+OW=$3 S_RK!*PDRX3UR7_-*%QD^G9*SIL 
@.,-LCBH1HBT^J+T#>YY6UWMF'@[ZUL;-$2TC8.4WRN4 
@B02!M]*0^3%+/>)Z!7O=^U]N$^$B3F92P\>NAVJ^,S0 
@Z77%:B61QV\6G!OT?X"I[AM-<LUQRO?;<.<O!.LP7-4 
@_S+:UW!Q7DU*WS9;!\#L,K=ZMTM@-WQS5;627)!!4?@ 
@W/ZCD*32E/X:!<#L>C^?[;>"@^/FZ))#@:ETXT!30.0 
@#9\2.#H-&>4IE@PBIJL+KC6<[/PH@N4>D\>;L*NUYZ0 
@"X6.%[,*E:/W$&:KE@JBV$88\2KZ(18%9D9\."/50'4 
@.-'D)\%3'&_;63#A3ZMGR2PRI02N4!R!I'T&-(UV^XD 
@[7(=\ "V6!=4:XA?IIM*D+U31Z1E]W!NR%@;;I5"2"8 
@1QN2^NN+>107IM0B$5@<1.T#C %-6#&87;^H]U)/\[8 
@G?TD45U2,OUMG$!2F47A!^3JPMOQ'T%AXYL_K:-1@PT 
@",W-F[<7589%9795'3KZ,\5V!$2E?Q5@L$/BHJ%BFD@ 
@)4&H",ZI0HV7HIP,:M-)R_\YZ%VX2.C1$W/0PDCG*M8 
@7-\_I69C*DCNQ>?Q7$#J=/)9"-&TIY72AL.&8!$\WH@ 
@=T<\Q=-PFV\WQTJQ;>S9O4=KQ';!-.QAP*T8WTQ+U < 
@ *"78)[.ZQ-35TGNV*GK"HK"8PH,"#=Q\#"*?NUQJ=4 
@7K8 :78]5A60-9=;?\P&#:.R6H6(_XD*%9U3D"UTN@$ 
@9G[$ JPP>XH=TJ^^BJA=4F FU#F(O$=MG0%).</CM_( 
@<BSF\LU4#55OJ=,/,6Z%)0SJKF6,6+)!9.>1#+;>ZA0 
@+^E#RNC#,1.H+T#72.6=L<<^5S:UMVYY<P)2=J:=9E8 
@7M#%\,3(\ZQ]K +"">,J4/;ENH/^U@1<M\(?%T*IW8D 
@.8/7E(G\=:.:W[BI69NI%>,')@$L 0(^UMM>3&JKEBL 
@S_T1H XTPS(\MP1'Z,M ,5W!P8(A5.8$=#2L879>[Z@ 
@:4)1]O'/&G2JO;!$7_)&__B?%#QBNC$L.V0,JO00.BT 
@PLXIF$U/GA3EWO=:DZ#$I%#V%F]#/^*2#/Y *JVA'\  
@4GOD[X)()SZ.-(&^^+J6V?9.=GQP+V\4T'I1IS@VT?X 
@'0L?4]Z.F/$_4\1B42:5BRMX>,2J.6V-5NDUGN!DQ3D 
@GLA&B"LW*XN&&B4O1;R1ME%#<"C7$<F#O^]F??L%;9< 
@:A%[F8,&6?EH I&ZOZDE%BGXP.@"@X0Z)H_87=)BAT< 
@6K!8-^D07I?;$X%YGAO^?MB&@/77:>[Q\?VOE]4G>AH 
@E#-]%$RM)'P]5*:H9,C(@T<EA-GQ1O=0,*2S6+6>BA, 
@X89R6?M3A7XZ;KLK_:,K*E7GHN9B5;?!4'/L ?FDVE0 
@F*8;'^W; T*CMNX:6ZR;TNR3Z=U>JRXPR\/*GFPO(M< 
@N0)Q("++EIC--SN/6H.;$'J% )EJ/%MCY9\ATT5$(2\ 
@%)RB=KML2[H(/&G-[S<01^1J/[T/+BU?8NMB0H/=;18 
@GWX<&82X\^LY6/N9[>=G:FGHS2OKL(@UR#TMD2K* 1\ 
@EP>IR&JIM-!NY9KZX<K$97_B5:"6]H32UTUAG_1E-,X 
@=\&BXVEP-@7MU4TQ,),;7YY4LZOF._G_F8 ^#:JXOZ< 
@9B'SB*8A](!7X$@EXITEG^=<KH#):4\WGD;>A5AT/AH 
@**Q45,A!7_W7G?$-Q@;Z9*O=TJP2Q=,45#%/!Q1?VG\ 
@@D2$TTV6E3^-.C[O(;O38!P_#%?$>C)NLOU B,<!61L 
@CMT3'^7HK'/N/VACU-DLNL8LK;)4? +D'S<L!,70]&< 
@F B;0RTXGG7A+Q;K<'E(BD#4\X3-#@SN7+X(?$4IMQ< 
@E6+FI-%_W4<Y>OH,SOHWN",\D154"RE8+<CWI,]: X$ 
@Z;I5*U<B0.%^?7'O]2!_1#G:Y+V81\(J;9Q#IRRFNA  
@I$*I^W4N HY_G:#*WNS^$NM!N?-I/(%LY:\7'WQ>$,P 
@D$7CWJ2QC84<4!:^:^BJ3-DPJ@BBQR!$BUS.>0> ^*0 
@YEDC@HUW]W3AV"CS@L4>:)2[=Y$DF<1:T3F^(P$UOF  
@42L/13]RO:D"OM*;OO=H%1(46(X9>^9B#_%20OQC9*  
@Z"26XP' ^.(#$+AS0E]T%@;3VU98.XVF*=WA@@A6^+T 
@5QCR,VMD""-$@5#+C'*C\UU_1WY!!=C=]U<BWU&-75  
@,?X WYNS(_LRDJ,!GX@[CS:II#/K_A#Z5JEKVR42R2T 
@0F]J9SPEVT>WME4(B6]%6SJHL'V>Q"ITJ5,/80^4%0X 
@, V*7/<;K#!N/+\Q]_D_7Y9J0XT>RNP!=+YW5(XIR2( 
@9\=6#W@4'-2C+B0J*/\K!ZDXD)OV3!7GSGS=!YRDXE4 
@#+IS->2/B'72MN\<"N/[@U?TQIB)UJ;H+-TN!2)DS[P 
@E2W5[-V2  +IR=5N0#)W4K#4<]X_)%S#3_G.EQ*&^@4 
@^A3O/+'>SL&1Z>)8W;%])O_H()WN(YRR1##2A0%0=V@ 
@R_Z_-N]I3P5[H2#;\'@%])=/$_0P<Z'6[Z+#^JHQ"]H 
@V.H;"[O?L_\]1J;C=D4D+ZK<-H@4U1&UCV@RAD=YW/8 
@TZAJ>1@TK)Y6(\8N5UV5&N%3+0*9H1VW9U8D9/P^);@ 
@&'?8M,>,S+&JL6&;QR?UL@.U_5KL.U3\*;$HPRT<3<@ 
@JH;(J6W>J2PY9_V[XTQRU,7BKO IS?F6EC_X9/U]"_0 
@;EWB@(4H]F;OTN:OH"1CZ24F*TON8#RUY?)1+=)^O8< 
@?-4-8O:NDZ#<I"&^V]T@&SM@[Q,:E]^Z(+LPJ(%!>3D 
@R47/]+QPTH5]@2P].,DU532;MP$GGW3)[$ C^D5!O+@ 
@:*C@9:C /79"/4L%SQ^_F>-CD=+4X#B(:PPXVZH4LAH 
@J0*GC3!0E9H71:ROFVU$_^,=9= "002OD#DR1V->1TP 
@"0+V>-,"=%!?*[D?2=RP^Y(B;)?;UF#R3G06+G35)%@ 
@W+]1C(#_S>EO!D2$A)JA%LESW13<CGH\]U-9%-*/NCH 
@5!B=1"JK,9$ZK9<:X:CD?@^-&30.G"N(W<B\?VS HLD 
@&B_6Y*/I+/)D_PW_%=QQY= U(XL)'+2U+_5VH!64&)( 
@0NOT?,&U7VC XCZ.B%BRY[.(S;SHF!#8Z'87O],LZ6P 
@'7AZGZZ+?I][#2>%64=Z-C6!;>$)GVC/G/EW6;.&J,\ 
@V--ERG9>M0S32C._'^2Q";![8HUI&P?K@<BT!Z  68, 
@0L+2PCP]>N)A]+IDDA(W$(JHE+/R@JZF1:Z#R7A5KO0 
@+8-WC1)&&6VA1(:SM-M#H/"D'D>\SRL_]@H$N^Z$OI4 
@7EA,79ZKBE98/=.\$(=482@N'B*C>YG;-Q[Z''C,V,$ 
@4Q?]MGX:Z4%>A:.*[F>E&KW3**(Y=;E?PJ&=\99*,F\ 
@B$8Q,WJ1[H2)#F82-CV4BT+I<%%^$\%VLX"0BDN<G+D 
@M-,\);;77LDU#(7$[#PGS>#=,1=6&'1P2'43>:?R%$$ 
@A!25N#SU;0DRSVDW>^&F$$[#+W;$PR7W5@&,Y-Z>(=( 
@Y=>3?.?-2W7_Q.%Y?[MIM=#H"!5.4L_$1 ,H[85!@Y  
@NQVHUFN145M3UJ^28-: 7SM)W(Q*G8B4#\E:U'4 F>4 
@]+NJ&/L:[TN:AP!C^S&=A[*UO^MZO1-'RD;:JIK\K^D 
@(-U4[=GM2<[2Y0[U33UJ?^.A#]/V8..,AJ!@_3GX-9T 
@<"M/CZ )*W@'SZOJ__M/^<!AQ1WWS3?C-7T')>=Z3+0 
@$=PD;"Y - **C=-V.2,!'E-Y_QG@Z'\)ZHJ5Y_,J%EP 
@N+?!WRWP=1[\N._DJ.WOQ93'$JK!,@T&<F\+?-SK)B< 
@H[NVO:<6:D2#Q=]#\/AIRI$AF)C._+GBT"F-8"HXXB4 
@S2'6JE:L5K>RO*\4]H-Q'^_VNSK9&X[..[-O]E$]\;, 
@M2TP?[KE)',6BQ1<A!<7#"WC]6+\U/,.\6J[WF>",A\ 
@"4-5Z7?AU)ER)  !*GB/GZT,2$(Q$%E=4_1@D#8+1,@ 
@5T53"JW&%>/3"7!P5U^H#;P6?9C?#7Z8UDOIMHG3-7P 
@]?W*@/MT)..LZK<\9\;:]&8O<MYNZN=L2?G>I]16,SX 
@"JAXTIRC+:QX&#%A,B'^YO9H49FX*+W'U<HU7CJX_Q$ 
@*5N_8.C:@D"D0#GOE9![TG2-I :6:DY O!!Y,.2=YTX 
@E?SC(MARU>X/);P4QW<0=[[TMMW/F%U7(PH9\E/]<"( 
@6@MAL\UA?KCG9BI7H^+J/U ?['2($V)""81>DE,^,,$ 
@K4JIDW@8LY95&4FRO2RT"HM^P$0%X_#S$RI:"*L:Y"  
@PA246O! IU9!7R:3QIXIQQN>4-@?$/K=H,T]^J;<<\8 
@?U>Q5&S+%$#%#2=X4&OTYY28>TMI!W"<Q!&PL7'5:>P 
@F]/T4!N/_;7G#<0ANK*&((%':0:%G%H2[[1XS?VBT&, 
@H%@:XU?W<R]._G><SDX!+RS@=LIQ%?,^)^M]3^DXK48 
@]!]R*8%PVG#O/)+]'/*[_8 _%&I'JV.A Q+7]X^/]"T 
@?GN 8_>9O4%]]H0I=,]RL-6U/*Y6^>*\BE[3D0AN=RL 
@U,VM&I0)O^CI&LM<$_?BYK<#2L7:]T=9*Q)25MEQ+MD 
@V6*F+LV%[-\*_@94TNHKQUZEPK@:OT5'?!6D3HA"-#@ 
@:DIEZ$:*7'X7WR +4A" K?_T/)_V [P 9.3!#53EH8@ 
@-5=HB!'*B5CNZ\Y+N^$P<U68T>$L]<&<=$]!T@38IDL 
@9Q4V;C^I%J('5^)@1PUJ*L*4JLMR>'_9JHO(ZEKNP&  
@8K*5\_49J:SAX@4X40TTTRZP\+7*GC/;Q)8H":-5<;L 
@<L4S']*;A3"PK,^VZZWR/%'G_\%?#<W351-W0R23[RH 
@#V%]X.J1'J)8WP)3&#<RJ<YG5<\B "J^%9:)H3>$S!( 
@!!J[N]_/JW4Z&$HU [WNP8T42X=(L$;WJ"HK5WR>S\  
@8:^@1FXZ;IG49_JA'@7^:PV?OVG><N\L1))<$]@39,8 
@L'<>0,FT%505A0?Z9*A\?YEWH^BWPZAK'7BSI86B?FL 
@'(KA T5583Y2E(^6;$G\D>Q6@$>#0T,85$;#*$Y0Z1H 
@/FQ=S!&@Q_^HFS#47>UQY+)I8TR14&,& E:?^6EE)=, 
@EU%Z34P,?E-W4$4Q%=</$B#?L40I(G.3L&WESSC,>=L 
@B'K[H_\UR&[8BT>_T0K78;;\<,G/XW][0X\R/<BTBX$ 
@RD%AI)R*U-/;_&O@Q^YQZNE.PG2FJ@))]51,.=79 AX 
@?7C8OHRU74:HADO3EP&+MU=1;&*4%:=B$RBT9#>!*+H 
@&B6=.DXHRE2HILP)"+Z( 5]Y/)YN,K4=0%^K]8$:(Q  
@YLCPGRK9- CS41K:D6L;0*"P&5 "FI^]\;M)-'Y 7>4 
@O\E#?H[(80CR5D >[D:@ZNX3DKH5-5Z.U0-%V.6/@PX 
@SQPGE=\BKXL!D#NQ7@IT?Y:#0U'T?;"5Z^RA02TF4RT 
@%XU1*D_Q2\FY5W9^R[*#W9SY*B,<V <$T]J1!IZT(,, 
@T=8>^Z[/;Q@^GPPVTYS%V@P%625*3']]L*6=O/]1D9X 
@85865?$@OCI=\^E F$!3"5]7\HV1<.6/XFZ?BHP;P%$ 
@B)F;8B5MBZ$1(-VA9OIDH;2!WGWSPA"$R?<O(623OT( 
@"MM31,7,P># ;&7GM[1U(5R7^/")O)*.H?H![2]:%Y0 
@D.7K+$9Z+#R_4TJ!.T0UWKUE&SGAPR366>6^B%(8@/L 
@%?,37M%>@,-0+1&'%=D&^$==9(+54FG_Q*Z?X%0'B7  
@_^WG8<>M>_5 F5@XY$H5_(ON;7'?-LF37VK6W@O8\M0 
@C%K'MP8B;,C$G^\K@Y43T_A:2*80\=),%3/5#5Y_&E@ 
@2^[?%4-#LK0O@3@"G?P30Q:2X2"*]OU:8PU>L<Z>,/X 
@XK1(Q):H#5.RE%N)Q2H5Z;.+P]6\]^$2]T&)^<V&]ZT 
@F,(R@/@OKN[&?7["!C$X$2L@$$!1,D;>P[DVWBL"OW8 
@7L&=JJ2T=*Y/A/[/YW_Q1?KNG^E8Z;D!V I>9#\O(YD 
@$T<Q8I-0*3Y2*ATS$(&49<T%/0!1?VA//3Q=9\4MK,@ 
@T=;E)Q6(3.B 5N7OU:6\Y9]U]$O4EQN(">0_GCHPTWH 
@47O8KI[)4:N_@GGW2P&M!36F<DY<A4!96:>IF&D$!UT 
@183AQS@;';WIJAFW*6%?HIQ@CX,,@"('#LJ##<1_&%X 
@$N%^SKUNI0Q2Y55I!J.E3^GQ&,3JE+T @GC0B*N^/CX 
@(LAI^9#)4JEI1+?P4YS(#/&,Z_>EJ,,D"0<JS_OTRQ, 
@EF4IJ@,;N"<2@BM<>+&6\LSDU."XH^90[7J!+^I$&6, 
@83J/=.77B.V,R7 =L "(&:8RBNPXWH?C!=3TA&OE1W0 
@OD$Y, V(2H(%'#"!SO8(]"@DJ!&'Y(C]5 (__D=.&TT 
@+RSX8.EGU K.P)U2#LN.FO?C-B>I<+L.;\%>98NJMF( 
@]6<K,_D.Q*KJZ=_?ADIO'JK+>_SEG8E:& @G7B"6+L4 
@W58\L?EX4D4Q?A]]J-S=3LHT&QU13W8:H_&+Q6JF0S4 
@_T@/*A6>0UN99*A[\UXHXUD5 +3JSB#YJWH[7$4'-Q, 
@Q6%KSRII%<#VT:<^)J[E58QO,QV*J.T%]:M2W4IC@5H 
@[\I8<G9RIXJ#W:RNSJ';135B.>7+GZ'.MLHYU8%'G-@ 
@RBGQXQWO,I8D"Z*@ +FCVG&()&^4#_PJ(5OYG0-P,?  
@1?1:=ENP@B$P\]VK&?9YD5@82PG@7^Y_U^L:%ZII[0< 
@5Z8UA&R"N+,UFD-Q5:GZ2^\2M3@5DE[&HW\@#H2;G9$ 
@2WO^^\MK7*QU '"8M5\RI/4 ;*D4N#^+3G-NDE!]'$  
@0Q93V*L9Z>?E5'M1'<:)LTHU=S2W=%P(MCG_0&S2K4D 
@NB4<O$W\\%EZE'!N]Q$IVAMF(.B(JUN:'2Z@^AYYJ-L 
@#H>0H^#WC?7[LSL (M(>"658?+LX!/Q2F<?:U*$<B/4 
@#5MB$'Z?4U5XG=!*DFMW7>.94R1]!HV+0D:Q6&KY5'@ 
@L\U5T*@4F"C^Z3GF"$Z]83*AU2G5YBEV"C6$A]4:G7$ 
@[X0-&;C*OG%3?86_N(8GUO\A=(H=E3V?//B78H7VO!D 
@8_D[1(69Q\;3)N,7S4 !U+"5'UUYLG0S]N"&O#UJL^\ 
@"%/WZ4.A/%3]TN[B*^BN#/Y$5/=1_VD):4ILIX7F^/4 
@8GN%Q,JQA\MQR-!#^1_969!U]T"P!<R[RN.<3[4_<IP 
@81D7!QPE0IY\^<RK\_"I9P ^(?"$W13P_E\G= R"UD\ 
@H%Y@@1C+5O6RF<@7\CC:O?HQ4XU02N06![!>MXE@)?< 
@H^\D]-R+TSOW\P6\?I)3D[_0RW[G(]7NG6DUYQE$_X$ 
@>&K-+[/7C?GCA6)2E4[,[1TD,0C.YH@R2)C;5/5\S9L 
@2Z=T@@'W"W=LP$N?0J3\1,=H$\W+<BV8_F84", 44H  
@(H4'INX4(T">,)5N[5I3:+Q0HT_=DX<X.&13UYFI=1P 
@]^:V/*9U[F,5UX]W>/Y3L#KG:<%0.0<9,Q0!^..CYRT 
@;_28%O(WV31I(;1-"K(/E\)W.TJQS2UK6@XHD8QW#U( 
@'UJKO/&S!=MQ[OR_E);Z@3&$LMJ]_50AW+<N =%ZWHL 
@RQ :@H+ACU"D9P\G0=F2X36 Q0_<D$Q=!T*3]!T&0R( 
@.^V>3  A"*M6=MM_E7=?:K9A?TPO+"Y>GI5^UZUW!=0 
@K&6;5,'@= Y>YAFB+T.6+"1ZB/K5&]* .+SF)L:JJ)$ 
@U"#TZ)<E5L_MZA=F;&'-+887*O.5.,AF#BOU]]PI;ST 
@JGAG-=7['<@JJ\*U]*JP5XI!2XJZ]3='G8P=F<[JLB< 
@V<()X'\+ZS(_GP-/ !CNGTV2/>M5]EYO!IY]K_AGG2L 
@X8X"8\ZH 5F'>*FO.^N"D:HSX2YE6%)FZ;#1/:(=6OL 
@34?13D);@LI@!!"C0^<.FUP"<];M*;B:/]^_C[*U9#( 
@)-?445G(Z&O$?4U\.)Y,O6JAQX'H)*0]TH* VI8$38( 
@UP[44LL/OK3ZZ(!XJM6=*1NC67A!0NJ'+#:&E%7JS)T 
@:T Y8[#(2J[G0_#-DNC^@L2@6#\2D<:GO^O>,=U7#ID 
@=MQ4!_CL_N$2D:SHZH+FXB]CSD<,MGI+GW@(&,:$7?0 
@,(@&5D?>.55Z%L#PO97X$QH8BT;VI4IY@,@>J_10=H8 
@61)@2N;?1**:OF1%Z5!N.0M+*M4VI*Z"MJ'13WN<)#( 
@ [^#7]]\4EZ=ZVNO.W\U_L*G[LB=<[C+I2P'0:S7--@ 
@$:B>#%4G/SF/Y5ZMYB. /%+=REKE"6N7S2WO/!%+N6\ 
@G[IF$G/]V03U/3]_NN"'"S87L_/0SHXO*"U'WPXCRR8 
@+](I2AR8:U^3L6S^P7X=]>.\%(ST06'3"A\G$:P\0G\ 
@)D?A6_7#;NRHR,&(K1RF6F@-]O'&:.KUXP_L,CLC/FL 
@M YOXD\3X>NZTCKA@.GQ6='!'V06L#WKG%+Z=_S*-"T 
@;# \I9+53=G/(/*-#MLE"YTVESKTQ]@TEJ81_UT6,V< 
@R_%?-Z5DTXD(P2(8<7;2&"(DVO;%?U(R#SOE_/_FD%\ 
@Y!)Y/<ZS@:/&,)5Y1 ,D0^S5JB]I4K(4B<\DQ(]JHNL 
@$/B^5)\.3T44 CS1R/- UZLWPXAQAR*Y[[$70>I+EB\ 
@6WB54_;\428^=6L]"XSU\;E?.WW8['C(FRNR\Y+DX4  
@_%G3TMH++_9=_)[G>$HDKB-N/[+)&8"A6]P4I$!YXR( 
@#^V;1FD*/RI-I^H9\F*QP@)W3OG*,NJ:[J^*W!<Q^2, 
@37)W7F!%"R/V;]0&'G)NC9=6;M'(I/*XKO"N3VCO1.  
@J@<0;J;#B&0Y0<BYWEGP=P>;"XSZEX$![%ME=%S4.+0 
@JLM6,R6;(O^_O(9M3OGX3VJ0N!D'@[Q+I_ , X+9"T$ 
@V^L33<:0SL^7AE2A59P@XO\#?!_<IT[#/&^;;*ZR&0D 
@]!1=H:>);DS%S0%0!2^VIMQ6Q*2"J'!+N*H)R"![_/, 
@:^_0%4@BHC4#ZA?NA#* 04M]O@)C80V[ONA1%P+T@4< 
@=8NM-"H.!;I@/*@]Q.>+2Y_T9O^&.0Z_!'$DH0;)%DT 
@G9B*V&VJ> *[S2&HL/?9>=4BR3)B"%+^AT-@?&Q4GJ  
@2>?$3;6,>F!;&+S$0D[DW;O+Z?2[--P#K\EN;7+ 2WH 
@4<7Q7.H-@1BFD&R=U]CKS(EI#< UY\0GU=4*9@*]0#$ 
@FLW6,\)-'-=UT*W,7L([98II5'WH(6QS?3YC4NF+'TH 
@BF=K HD7:;>(XL)!9+:5A#9*'9(TT(ZF2X%.;G 08., 
@.'4#ZZ#$[(I20.,G47X$'$1V\U*HN<IQEC'1DY0]42T 
@VSPF?99M[B5:40Y\4']+X)H[GI5Q?TE+9!5%TK&IY2@ 
@E[N6/LK.</*-^?/KA7$ YB,W$D?;%4>RL;V .6QGMH0 
@!L>?RI W<$KQ-R*1[3&?5#%.?3;X<APQDC.O 2%9D=( 
@H" > "&]*%MBVZ["+T,C1'ME:C$!%#[(IC[PSO%KX/D 
@UKBK1J$79DV,7G'5!^#>@3OUE=M&;]>NP!U#\UHM;C8 
@[W[65O CG^6U_26=22!Q$M+(@ZRAUZRO\]UTA3FV$,, 
@2@C]6P:F%T%9AD>>K?1ZD8<7&"P.2,D&G>F!_/YH6ED 
@CC8G8["V&FSA:4AUL5YNX)MKQKE"T5M[-'X]Y35?]^\ 
@J2BR,@INV7A"_; T%S/V(( ME$[3#.0E/$G8[:=:>1T 
@@)(*4K-=&*(@;*#;#^ZMJ[6ZOWO%TA7#PYENQKU?"X0 
@/QBS63IC"K \1%*MWD<1*:*;#3)<-UB*V*TM,?C]X(T 
@=D(CT<)R?ND7)*\"U0=XE*BD!"B:RA?EJ?Y?ZC)RRF  
@2WM6X4L :WKN)% UHC)YN! -_;STK?X+23'5J?+9KN\ 
@.\2BV'?;]2ORM^HH((-82,IRH5V[A]!\JF]\SUC4^UH 
@TCAHK/+W&KAZ(10=QK( ,L7A$(R'=,JRO9 9*]W+!RP 
@O2Q\O]@P&BKC?=/S-19(8+H+JFY$H(::$AC+NBD'4#L 
@R5YNVA,$Q4?67*Z4NP<2B6R&X"^EV"=SU6I3[:VSM<0 
@L#!#4E6S'WR_36^7XI;W(=@JZ$AX]KJG!$ 1.*/P.PD 
@$$'+43=N(K\^/RP0A_3AZ.9@&VY!DN#PB^]*\&3<CA\ 
@#-C4UFC:Z;!$B(@9V3 -/Q>5IM-,H6!_&"]V:A5<MMT 
@E@90K!\'T^AI^.W:<%WLJA=Q=*HZT1@RN5D^,3>]Z\( 
@N/J 8UU$-@-%H+^#%UH A,;@^! >@9L@V'V\)!9(BE< 
@ZPT !8YLY$]B8CUQPOU;EP[M[[!+.030Z1+6!,Z \%, 
@WEHO51V>&W^HSVY/LT VPMV4\,TW? $J5XN.:M4@=?, 
@D"G'AZ:24TZ<%_*2R:HU==I1Y&9AZ-)80*0^RM"$ DH 
@-;A;.8^O@12Z]3: F/==,PROC.!*,15O?E*S"@M[[-  
@<4QI=Z>X^PMM? 3)"UQUY:A/M(MWSTEY0R7UR;BD7#< 
@#6PPMR]?<?^\U%Y0-'#[C 5#EK+YE5'%ICR;T[MTB[P 
@"M=*#SI]R2GI D^=-.3F9)5;V57&=5\%:+_%BC>[J#  
@*M&;V7I!A4V\PC2L!Y^.7-<3C-= !P'2)V<:])++20D 
@R0J5B2W>H]< N3%I<F("TU#&;%RF[E_&51?Q4S8ZY6L 
@7\&;-VIV#8,GYB5(G%:2-PB2"M&GMEF [[SW5^,[ &( 
@L/G&N.S?]L)S4=H;4M3;J%[)??01Y*-.WSMBIA;[FW4 
@9WM2$2@ B63FR0%QK0+Q8Z K Q:9R2O.J15(+"BG94H 
@F$=)#<2<ZL="^8.IH.M![AM^V "5S>P/=2(ORQ<-  @ 
@-UX\9Y=$!N+\F_<]J$X7PY5&03NV(O.C;6#M:GG/Y&0 
@L6(K74@, L4&\%>+7?$;G9.I>3KF!]%4)Z>U]%Z+?LT 
@@-X J&0G?%)( 0WHFRS)%N8U*);C@@2)H$_G&%\@.Q, 
@. %3RMXH1 %97:-]LX;T7JJDVZ]2&U$V\,AD#5++<0X 
@+H57@]A[DO.N<XF[>SC>\KG/2$P=+>KWXE7HJ#CJJ@X 
@5A7[I+6TB$LT"]@8M&D.XDVE(2JO9TT+WO(E'')]^6$ 
@6J15JLG1>L8DJLCVS 0V-"1AT\.'5^T$_HZSXE_")Y0 
@&2'*B'>X4\ =1FBH&U9SO%<V5H2PO>:*&QFFC\Q7D]< 
@BXL_=_NUUI028+DT_I'ZG;[RY:_FMP4$NN'\"#'SOGX 
@H$G9$+3X51/&H#$J'Z:AS%[]W\ Y^EK!J9ZIBM9)4K, 
@KFJE7X[CU!G724"7&*-T7N[.I5/_E]E^/':$4^UD[ID 
@^=,NV(= :$TVPG+B^.P+"9AA4'2XX^QCC>[]2P^-P?< 
@]*:E29-ZG6V4"E4V3QHE&TA#-,2[]G?<6)-2OE%%=X< 
@-6BJL'GT4Q$]JD>0EV96'RS*M<'0C#TOME[(KN-]9JL 
@,)12CD%,?63&<T4CT#!?8UT=&$DZ?E_>;AKV@Y41X/, 
@;26 2O%H\G>D*\I42K=C\RG8>+Y,LBR#,%I25SSG2G, 
@KS\MJB6!(:_'QZZ2 K(5TK+12.\NS923P;>W?[7<EF$ 
@![11I'JT"*J^*-6^.SGA&W7[ZQJXW3X%"V(\;T=YD-$ 
@<2N-HI$BJ1Q6^[ (6<ED>,<C6<YUQD^2P!9;!^W*$/D 
@^&#LI#]QF,[S5OV?>WH5V'GJIG3%))0P;'=7#*">ZGH 
@=)RL:I"SNL"TO"_'N%?=GH+(;:-NJ5R9FY@)+#.$1H0 
@:RO!G%C#)XO#M5S<5C-A;MB\N(NFN-T3V\='#.SL5!$ 
@O"VBGJ;\[S/+G=J&,!67PUN0D>BFN@P)\5&%RK@/]!P 
@'8!!3;[S5/)YUZ:JG7OC@DJ;!F @B5@FH]< L)[]F$0 
@CG5CU:BGM$8&-&U3BC.B[ X7 ] 73$+>88ELN^&)!"L 
@B69(N<>=BP?%(X/RIJB>1.$]G07G)YX) 9 3!F]NE%@ 
@;GB2)+87+[RRSL=7)E.'$\[=@\W"&+9&TJ;.(^9G6#\ 
@17/F8Y6Q0X$ANY_"Y@2!S@=(MN4D;KX,+<WBT5H5?:D 
@6HMQPB#Q-JZ(5K2+J8RB7EFG]G!OU@'M?)=J!L%3F$X 
@L\+KX%X9[%.\B([W/NG,\L'AA8X6Y/!):%.1O[G)LW0 
@^YN#V^@W7G;&IT127 .;O3F52ZT",TQP\-P-E>[77%D 
@V!,DK-)V!*)^V^=@TRND(!&^+CL*L*B&*  _)90-W,D 
@_0TVA#&[U59I*RN&+E[>SS>5T]=V"U4'T$]9C ?12*0 
@-;7 0K=,799=BS,K_+WC1I0BPOI#5)Q/(==<3A@2<;T 
@*8C%A"><(87O<M8Q</GG%N=<N594.+ZG8W?CA.1>G,\ 
@5=VZRT\9O\D7Q;H9ZI;@4C*"QI5?I%T8RIKGJ4O574H 
@,&3&+[:TC4M:'K-F[ODPW/7N/ZB5]+_/:CTJ= -/I6\ 
@OGQYC_04;[,8-*<Y"P_<\UX"^P&"M._R:S>=JGC0.#\ 
@*B" 4K-I7/XFF!ECQ[@M!]"-/>&\@%"GGZ+"/PY%W_, 
@O@GR](0G% !7[Z12)9O:V@X6/A].KTY%@T1@P(Z(KI8 
@%._]&P =5[8=<F0(@4O<8M_ ZFW>KF:)Q1]V>W5^E2P 
@L=^*VT0\T$SMYU8HI0.TD9&,,1C-YSX3I8L\7CZPK_\ 
@?L[GC-? S7E1E<N*X_C:,Q8R21OC!FZTUXR!\&1L^S( 
@(?C7\,3R(DQ=AB7;@OL,,%EX'IJ .8"%9/Y0N.>1W70 
@RD[6@NHV FT X=D?$C#YJG1.66(2'&^/G,LLQ.P)'>, 
@@I1>.1_! )=J,Z9LG-J]TZLPR/*_(D_]J: /91ZB9!T 
@D^\V-./J KM@-([:+M#+5SPO\6?<FH_..3Z>S(>094H 
@1_EG=A@? A 'GL@D+=70HQNC3T0.U;9):[DX\E5M@%8 
@/([0\9G.JD6K@D=P-KY*%Q]TV8VD<]=6D05YPMRWD4, 
@S5#@>K0.-7OCTKB-D#2(6VC"-.J@':GZ>-8\+&580]< 
@/*T57JOX<\!+;+<&.F:Q]L35KR\/VGP6O[6HC8$;1$$ 
@KDU'+I&Z1D#\)9M3)THO(LA9,BFG:J_>0MRN>L-.R<4 
@O'4GGM@ EMK/4HE+O& R9Y\/AC]@2"F"Q<!4_ <9+2D 
@[.LK'=8A+!\ R<M6BPBU<'%+)"2%((&!8\X II5%M[P 
@6EM8-:]$WEP.Y2AS8I/UXLSF.R<FS'TA*O@]?BTFP9H 
@JJ<;[M2I#N4:,*MC2&6'X//M)(B Z18[/J8QBX%NG;$ 
@5OY'8D].)Y"RTRN;%IW+E3U89H,N=O/#WFD-M1A(8%@ 
@ZKT$B@(-85S)2YZNZG(G /MPN$9,+W"G-F!(T16_Y>X 
@-9]?MK6H;U^+X"Z-B)/'"-C]E^(5:/UEV>C0ZN"HN'@ 
@,]#M/YEBWWD^Y[JT&/M241D()1V%67)GKB3,S"<I)0\ 
@)GVGKW-6@E-WF.<0$;$2/@L!3>^SZNZ!HU%9$J47@"4 
@DJ\C,9#V%1A-V5SMC_^<>@ TA@DA68W%*-WT=H=DSW( 
@WWLQ.:]7Q+)(Q;R^I,VBVF4D#(","MKH@L.-B8Z2V3L 
@Z6C:+_V!1[G(\$OCC'LUV5^+2)W7D\UA-B6+*'_(V08 
@:KCL(@;^FR!S9!(HR-C6'V!^=1'?I[N!.)Q2>2-$8:H 
@)K81V(/W*%4V92X(22:]!C6I9K0"KE%^P:B1G./874D 
@6;N4)YFU%%Y5TN'EE[R>#W8,^,V&7YF80184XW_WEG@ 
@OIW"$"I4DB,0.N>W6<043+?1!:[CTL#)KO!&F:^_D $ 
@ ]IVE^]Y,&M/_&\-%@I&Z_YD_.\D--XO_0"0)?OM*P( 
@(9H-P6:31NQ9BDOM:28&Q@W>DI,<!'B0==%-7:K.[_4 
@%<2K5/C&Z'J'"8.22P %ZCA /4>0+NJ-CO:&-L]VWI@ 
0G$ZJ65<+U.;'LWA_ MW<S@  
0[?V6"UB/F^;__1(Z _+&,@  
`pragma protect end_protected
