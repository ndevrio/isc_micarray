// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Sun Sep 22 20:49:28 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RgorJK+nGMhghd7MaoVdPy5KDUdvucFXLiVD5Qw15QXme+NZx7Vos0+Zc6U5txAI
YVx6TXtQ2rYhJYoEO6pvhyLTQ7U5L14mPRh4JNgvDPmTiHXd3XRB6BRhCTB3/Get
d/120+1SBl0jwSMLe5dNHwv/d0i/kn5IcIBN6P7QQp0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2944)
xy41Czp4SeOWWKVdYLyMwpfJ+lD1hkMHEdPVNIFTBpnXeSeM5AgImWXG2ixEhX1N
LkHb++GOiA670TzsIyoxy16FTVA90RDalivL0wn0LGlX7m3mFPXf8aN/+cvdUe6d
UF0BNT1tYUJZvjpsnvPhxsFtgBnepg9k7hxd5mr23XA5byVFaWAOYuaJ5cm0RAZY
4MGfy3yYUCg2+cfLZqo5Vr6HnAPCMzbSe+AzBv2SqPByxGHiSQmmpmz3/H1yQGXI
D4LuUgg8Kjrl115pNgJfvCMIs+NzUwd0m/2474na6ZV5gIDpwHOJj7b/ZHloQMC7
d4MTMGaAoZTr3tZHC/kNpJUdMujCJo3YVh7/Lp1hVUBuDeZO2P1RHl80+AyvlEoQ
wCKDe32nVQ1jTT0MNPr1J1fj6C9yogCwtF2JxedBJd7RQkMgqgGizoypeczkUHR9
gldElDubamgWCAOfIBqyESZccyV22IdfR8qL2ayB9jgkz7Qm+Emp/bH825CSR3/G
6lbSWFkrlfUjuiuHv1ToOYYezZcVxWlP8COtSZKefib/ndpZvJNkGWl3yndruNGB
FzWak077bUFfJ9NVTSMOpV8GQGI+7wuwZ/Y423NY7T2TadXcgESWbgE0m2gNIPPb
BXLwNPMm3CDQHy1rAs7Cb3mPaoAxhJ93I65NQnmaGyZrixEmV1cYJXFyHT6kp0u0
CfrxHfmLxI92D2gVYgqkJhDHqCNYPLzD9VxEXUuG4w6GGtz/mo+Xal9DYPhG747/
FjPMhSorRv0hYG6Ac8+mH12N6AJ2joGxTz/HoZPGhxZjYMdDfAyFtuwSwxch9yuU
NQIcoqX0f3vh9NCnp4s6lnc9Wch4Ar6g7g5jwvnwNn/WQrl0/3pNF6U/aiJG4rKq
yQFp13dqorL2CShVHTLJlYNMfXrpmq9Hk2RwYX7/tSA6kFSa/yb1bl+U/Ex0lqCF
V+Yg2o5bsn/BU79mofSY0nYNsHP/wLko+pJ/E2FqjTQ5+qGSQkIKQ+3ZmEiMTFgr
4LSVbJRnBq27iNUkKTJ/zZMikAE5QSFwFncz25V9jko+6jwsGq6Hck8CvWTM4bST
2FxfwDyO/eZlGByuR22uS/xXHNnZLz5erbS1XzUYqZ+WalmS03NJeQp/5U7Mqeox
0Bpq2U35ONMHui6069h7HL6vH7wN3HEhfoNFnzy9Psnakn/iIm4eDkYYfiAAM4e+
vCNx8BOuQBVsTy0NiAZviCz0t3k1jqDx9DVLYObu/A/amfuUvzhl+oAvhDEi5uDf
steqP+rFmOuzTR3yzGU4mCZBij0bQdZ9mVgrNmEbx2RcWpBVvbQIqsMvae7pdpce
ablXqvSCV/EU/Ts4nUi1x709DoyjYn1nZT4+yr73LIVasGUu/RhlbDuU6rVnGJcK
/6yMtunFtMaBBwHpWG9Dj86Qu0mfAeJvDMDzQSepUxHS3Ff97l6O+AEX1M3Q4zvQ
n8TNy2IFFB0uvVW3EGaikwyrQGOzJrlW7jn+xPFm4sNh80iHEgICvwJbSQOcFWS/
GrEam0tLXKb4IJ15eFKKRgE+NhiQ3Z/efROpcC47/ewnJdiS9ovcaLK81spbhG9t
2urz45EpOCpzmIZugpOJiwDfz5fg+cDrfVSxcGddFL2tqkzEA4ZGFx65K/1O9m9r
tn0+z1gse9DQyy4i61cgmlkVnKgR2oC7vQzYDZ9TwMb4t+VHVr1m0haWPyHzSelt
9nlY17e9W66tTBbdxYEf8foa/Ro2D5L0Oc/eH/DbH0ficQ4zbarE0ieM3eRtB4cG
O4BwgvD+yV0L5jrIZ0d/jiMAb7NP9/74KE/dM/vTV1uzQT+8gmHy821nqEuH7I07
oH3SQ5O/VGUewvB82iu12r3Dz/+7QohFIB5BhJoR4WrFHMXtz9+no1zycmGIu4DB
Q0Z3z/bEp7TIDfDiQbr5nvcGLXO20fsW08ciDWiPYAKv/UV+RIwUX4+OySCCYUqO
2Q9tTERscnVR9xWhLo3uo6mC8euyyfQHhdq/slNGTpN8ypz4DwErHJjS65qXAPSv
1jBT111DSVYXrT4r3N4CvrYN8lMOQpAqxTiypr7plkqsxxc13oO7T3FmRFu2rPuk
EGIAu+wEpkN53In1i+QBkSWhmlKkdwWDWhf7RrhtP2PVqUsayPHJskBP5fnNzh9l
hwjH6hAOOh8kD+FTQr/jiH+tbWSsTINfhQDAePeCdoMdhRF5tQymfiZMNu+Hu+ij
GHOlDW/vs0yeuvxaC//CnhYgW1RxyW3kU3VO+eg5wOKerHWmiDh1t/ZL3VTiGHqw
7ZXQbsIY/8RBsjQFKB2j8NchWEQJ56TGOXSzjSywJ3+YUNoh4VdPcMzf7HgLiXZU
bzzc33HgsJcryaFdEu0C+IT6eCVXmVCnkOdyFibkbdKn28wXrPK813RKCWJ3Snpm
6HduhPVX2wro9CVgNKTN1XM2Z1bx/C2LeoUy56Wl8d7WdtaipEEk5gv0Cxio3C/7
BZyrbFgYbDmrEfTuB/xtaXoOINWLSFSKlmXq0/r4kppoKETbJI59dII089klj5qm
6Zoe8aTaEDQbXvMBlu4P50SECHp03LuuxQAeUh767W4wNtoHfShkzQRYspGiqPtS
6q/onF18zFOPUA9hDo3D9Qsj7eGop4Bix/gL5gYXZOyRf6MOHrpv2HUDK8/Xw0SR
Q9MbA8ZtM3N1AmRY4POoknCNQL2zYP6OZFtU/WVyDs1Kk85i17K7h2i8qwyRIt3w
kjxZSDUZxGlcjSS4FVBqAMPpnSAXLJ9rPPECABduO6ctezY24c7V6TXVDKUXOOWD
txC46G59gfTZEZBjYytr/fH7MxlGcd1Mo842HX8MBJPbGssP+1Pcf7l3sJsHs48T
rc9VCQuqwG8oZYIrIBjGRgEMpBNfrcQP+1A7y/JYrc10dEseyR8uR4zLZM2LYBw9
0EXvPVVurJkgWj642nGjtVnjLefDMR9+NWmpWFTW32aHD6TX3mFdro6x4RHKjQtD
S1FQlzZSgqRnEmVZRVGxekmbqduIto9rOALoTAfrWVBskMlFwkk7jk9VREyIwNQ6
cc/5RjSB/PmHXndmYk7PpSCOLjUz17lk8u9160PPoD/D+MvGUi9wU+erobdP9xR9
YXGMehIxwj9ojwqjjjAccSQZgeT/dQf9G/ljPr8vOQOPmlfwaRZNL1vM015mkz5D
FYAg1SHjvdxgcFPy7ZroxZNvEHTcT2BEkCic4q/Ipq7KKlyg3ZjmNqE35XrS3tyo
RgsL4vUwmoLi+wLts5Yo6YKWuN8xByJ3XH3PLu0oB2t1WKWnXeXA6to87zMfSs1T
qo6JAYXeJuW+Fftnhb4ffXH5yYhmeFJNcp1X8TQew9U6QlBa7OPXkNqhjtZ4Khr5
Na5vvddrM+TSte33pvWrjaX5WtG3CGoxkzLmOhAjPzBjYv/jgfHKiu6LHV5Dr8JL
fhtFr4EsdWH0WvT5RYZDvDA4g6Ogf7m4uPrBaB7w9xyDbF2RNdUALkVar7eL44nk
0QHKdjCK8eJf2TXmaBvSzRT5WjFAuRjudBX/9SS8ks7CfnJ3//DeVo6cPaLFIQ/S
IbBy/jMZvkEPmnotFeh2PYAWlLSFGy6T+bcehH6ZFW9w9R9nW0rSl+s4sJ5sWoY6
MLEZvBpDxVrg1CpDcTX5+ZrYi1yfOBliFGHRXt9DRHOcn2NRIo8BFC+qdalaodys
kimH2aSZkzm3Pzr/KQ6X9MB2rogvWcGXPfhQmT3smeldqVw1nlQwv1p/j3WCSikt
7v/aULKwNIZ2I9fk2KiSuUvV/VC+K1/ruOOaxEctsI7nQ8KwpI4A//mylg354VZy
yHchrl7Uo2RSp4fVD8C+fJOWLeorXzKFaY57GrcNwgSe+UXAPIGMt84JL5GxXYMF
MRoJGsrP680vBQe5cuMUpw==
`pragma protect end_protected
