// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Sun Sep 22 20:49:28 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iD93N7XDy5DehzLBAvjCHn45I7JVG6QcQGfDQoRxxkTZOVZ45HEasQNOEPk0jEhk
aQNpSM6YPAGsFWtIU8cCQNMazbVByWQJUH3s0oULD/vZ4ubtcgHnL/pPMVsXU0Aj
VtXDgASL1n+drdq4G8DzK62hWFwVlJ+lpAOSznPSRwg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3008)
YhAiDWp9Erv2TAzB7pKQ07X3FOOMUOkRjUePcE1uceHvInFiyYHMVHAy7e9w7Nw2
bcRVzVhABsHFrd8/PCU4XqLUXyIkBncYBRzRQ4owLUdO7vorZLfeGuyUtT5Rb8YZ
3f6eUSQIYEaurWWDRcx5PMv/44XGPJnnwdN2LD9O4Rl28VQlewyUyYViqLIGOoUp
iWUyQLWuHrkDUDYRpHa/0bYYgJMxfuQ51D34fp6mQ16qSyC+VagEyw+DN2RBInB5
3XbVx29ZRH/zKAMsBHBJ/NPWI2ovDKlyNdD/kxlxX5qzQ1gbxTct33pX9EoyFHBl
a16YC0umChTdlF1P/nQ8BR0DRC0HvdzipmWcl6VblYQry2zTswF5rR3K+LzJWTvZ
q8KIuckoE0cjFhU+SaDTPg4YHBwwoR6j9rbVoQLBdclwPO+PZ8F7/WW5s6NvdjU8
X5QpOmHqqDF+iq9UuNXIN0ndMyGbCHWWmkH2ujaRT0Z1hIFX36UyaZOWSVcp/GwR
Xqj1fvQEq/1ol4zIoth3Kf6HxrPEsT1DVuEPnZnqPK2Gcl6jhbtHzouxiLZ9PON7
GZZVL87aQ6xskqqUvO1NKCkgu1MxvrEUggZPoq9RYwalyLG5I5NbgzQK7IJ+718C
rhp+FH8jqWApk7dZoNib7FiAg8GYIToOoRpLiUuGq8RxsYh56B4FVYX5kpt0yhM+
bOQ/9KQWNIkzzCp+i+3fjiUkogTuA/h8TSQzCbOX8Hh3k4bxsrnbpc/O7pV1fJ0r
haRzKIqsfp9cNeJHPbSk6vNaDGWN9KzeZi4VJOCyb+QXP/TMGcSORagBosgJDef9
v4JZbDGzYbRlWA9fzGzPz4Rfg7nHuKKwrgdC3F1u/mKYmDmGlF8NK9iZ47ImWg9h
1uULq47ph2ui5YglnJ+csNKAmObjLHGwJUCTuqydDasz0z0sDvTT7btxytHnI0kl
/y5hldtEGKomoCLgW64Hd62oYlY+TSTO0LmRl3p1loLItEhxl9CFMN6jes/PLZeu
1a2pwvLvWPYeL6yJOefzn3BgT/xhcWUKIwn+FKOeHBHwK70ulQ2SlDS+nZ+uRSbI
3VCvqRObln2DZWlwfaSvakhmzGEbaYZgwsuw4ey7SuaMtc+xR5umedM3ygUsm5a3
p6AKEIw3JfPBxrRjfo3MCcRJKO72lEH9Iv5CIgYFoDYYkqDi4suFSgRPgtBUB0Jj
ga3TsF5+2jZuK3pqVNpyvlj6PgSfNQyymI58LmmnqNB0nWAm3BTf/BkZvHJ/Zvf+
Ps5geFNM6hMdjY1JGxk5nU1/4KiTEQiqUJ3p8GF4RCuc8d2Q38LK5jCFjeTCmzb/
V9Db8oRiqsp3uvaC5SWt1W3+cke/RqASdeBC580gz/iaAMJ1hc+H2Rt0HzRoirpJ
T2C7FV8z3UkK1lAPQOCnpjz2ow2h98vjnEcBT4cHQdDtonIzgtBsStCdjTHXxnlN
BHiqg0GrKMifPRDeeRsgjNd/HiXQ+b44/WT/qi8WuIyE1JWRImxRi/Qy/LErdP6q
iLHRUrWyGKcyQyNMSp+v4xkPh5jszmpguD9O4tm59Nfl0N8C2RvqJO/cKOMFgzVO
ZltZjttSZu3sIT5ec1K76dBsLw1ArvpBTnDqTpsHiaMp3ULN1YcI07OLbP3BmDRb
VmE44w+kE3mxFlLVVc2LqQNwzWVwXmLE8hdIB4EzMaiMCYV1hUSXzoKta7UVm0su
2VkZjkWZsnL1K9ZFswgByxApb2IMYo78Cm7YUH2lF8s5ZSW3vR49HT7Lm1rdnqom
Rue5XAMHLJJS/OdDyf/jFUvZbfbL5qZ13BXNq8sfwK6hJNjw13jdDfQzJU5MdmUP
AAeInmZbKreVqwSiLq7LTPLtBdUXXzYZKkbECOwSQvAbKvAsH/RHXPYREXgvE3XT
4mUhGPG7KeLimOiOO0rxk0dQb1Z8Ve2AoWyxvqHq6S0OPO27E9wAIRqFXtrmB26t
2nU6LDOoMCU8WXjSoBU3Y9R954YfP2OrPopOcJhbHqdrNSnC4cnwYevQ0zE7cWwW
/uOf1Bs8e0b0I5PdZwXA+d07EypcHzLGsu8Wb7BLceHco+TjAY+ny2P66yJApZKo
WlieXcSnYSoz7Nfhs21H6ocz720GF6mhbXZ2CYtVeEaWJ23vJUxBLvVIzVYT6BVT
Pr6206AW58FNZ9D9BiMqF4toH3YdQTeqg2ygATw+QcNno9SIVGlTUi3wbBHcAEaU
md3P5DLE0VaBF1kNktdH1ZOG9/kfrlPMJrhQknk22oEDCM07ro0uTZvHecDa4emM
9ZBSDCfGBFtp73LVtA8pf8Mq7+rumi4IT4dKP+XpcTSLhlGe3Y1QF9JueueSD4dt
QX0DV+6a2XohrP72VdBxMh0jJCf85IAUWJ2Xh5bU9G/do3kQYO8IJIeZgV9esAw7
UcR7kJxAK23wlU2dACEEYNZcyL/bblIAah1HfSfzXflwnrk8HIuTzLXEue1OHdIE
t8B60dmdhRh2a4INYv0Ot6kP7mh16XmFWkG4KpUzi/vuanB8W/YQy7S5m9/YqoJ3
lwFJFvnO9W5x1AfuQ5rIH5nSXHPQy8o7maAdGJuc4P6Z11K7GvN/U8CRlk/WWjC1
1AdSXV0HJM+yMG0Dz0P1SvtP892iqFkHQTAocScm951b7YVeg4p38pQL2sLHGarz
v6fhgDtIBFiXmumH0wgY8aRFEqU+pg95GInF5I+F4edPXCyPMEW/QRG2FXs08OXz
FpKp+8F3F+XZogVlnOmhpxmZ1XPMfJaiWBGeZnGLXV/BN2J45veL9SMD/ilKFRRL
08Sr2HDpYFgWrn6ub3NOq4O0dblEFzKtT3iqC7l7C90G94++1fzF/kIJ8yd3FhqB
gmRiHl3apcZq1no0GSU50kjivHDafwcvjjkIazIXJHhhZthT9AiPxDelVKetbzDA
QB4T+m0mt5occ/two0bfn8cOj7y66uwhKT203CZZIwh45XSRlU0k9MVkgzS0yu+F
7X3iI8kcjCu/61/OIAhp+hzjFdjkgQgHjdyyELCNIYevcfG6yVMH8dUDmUdVKb8b
uYnvNzp/r8TcyARvOE0rLRSga+dRAz1s3FlVBtINEtKoYTmqUlrhx/IYG58zy/cM
2+BG7xhbD86GOFfvc5h8bDTRreUUEM2GTszILICvhJJfKg4LHJYgBJIzVrS9KE27
y524BTQxGsS7rYNx8JQ1agIrRODHL822ZSNlByg7KhDi6ui/+YkB+Fx8EqColAMy
dNT4Lu0KzDv0lFWnGONdqqFppWveMOUWzGnFjpYglyAO0cvl5lXz6bXmjqrviE0n
7nMNdl4KkanoSsOIBH4x4nDC41v5VhDGZaiICw4x4CEjMd2zhGl4IHhPzt2Rk0LM
PcdZ5OQmOxf94TEzsdUiyIppUiiFQXe/+ea8mOPa6u1/hKGdJH6Ft30yDETFUgVq
wk49RC8z2J8zxqKhF14fXxVU6S+hyo7Z02pnpt+zMksjpnlF4fn2u27x8Z7KQ9OV
12YI313bkbKaGfBCkSysm54QZ/yke5jK75m1ROMf6sFs43KLO9YGO5/PdGIFmCAl
8oD+rxS3X+MA667EJJixy78C6WUr6eZeVxgSvdpUgJq/5A0qHWjpN4Ezh77fp+/J
kDy+dUy8EUSFgGKApzVxIrSvhA7klNPwT07fwdCUmq7miWJdqJUmZ0w1s6hRe3k+
FdoLeww8yKpV7qSyGB0Q/hpaQSxa4SBUN1iQr36LGi2xRMrgjPnzfhvTKVIvQX8S
FwkEnKvimdqJo36OSfUzw6i9MQig0s6vUHO9IRQLMLIpcINPnCNrAy/diico3jJp
wRUX4YrXljhEkIfcqz5FyJVhR9T8hTyGhcZYV/MdCdyWFD8pqnuCAeieDqsJOWNU
P49ZKZzCsgAe9w2BE5pA+ITH61w2tC4RRNJWN5WUTmZnMhMymt6JtLB2WHhR03Q6
hSpkCwJWVhmHsa3ZjNNU3SPFEp/XKL2KOoYU3X5EMGc=
`pragma protect end_protected
