-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
nyJxA9CAUIhiZjpIwzaCd2yguhyYmDuQT0Zv7Zo3pKwrTP6jh2Ss3osAnF/56qVS
59M2ihQ5x/xcE/FZ5l+8uIy1PUg4UWj8d+yJf8K1+E1Ltjj2YE7yEfNQw+475jIt
M5UAh+bo0W/vD8l63xr3peIXl5y+Lvq8TzrIQP2akRc=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 7488)
`protect data_block
r2YMnjXRO6zxFO6d+16HG0Ssw3AxGgbzxqqHU0tSlZ3pZDsaEVQ7w1zgwjh3RY4a
agxpWljcXMgBDVs2rt1gFP+znM3qxG/s8eQ5KCw72Q6OpzLPDB5WGthJzO4yZ6rF
zyOnuMn1wY+FT3yJWIB9/m7qkaL+rAA23pmlA/GXqf/W3v+a0hfeudRb2x8tvV/V
rIBvxdoWMX849qYPimpHu0tCAkBYpWXYIxydWMpwyd5zHbqGoovSpKsJJipPtb3y
P7zdD4HZDPr+bzMetqlTdqEIZ1j8jIrb17PwU5mxEty4259NECNryf1AGdQB3mzD
fK7Vtl0A+AcCXzYX0vn2RO8Wm/fx/wZ9A5bNoDmYDqVFsY4F2pLuCcRHC1kGraMJ
FgwRPg4E/pI/7IM9JAnHbSKnmdVnvyh5iU25KErW5YeqxvfCza6JAgzgnOFnXKw1
g0nUZdHjdIM381cz4oULb+xll5DBO0cCuLEgNyAvPv3edkb812mSE/rZJvVTbGTR
KPEXKiU215yQQeUGtlFHJJWandB1HayeLWLWPf7HsDQeeNFrW9Etpt62CSNb+CIV
9viMLvOPf8UUAeVvQi8Jvr6ZxomRtjpSiSPxjU52qTWqyPZrWM/23dZ+cidRqxS5
dNtfeGq+oY+ZIQIauCCzRvpwi3FE6jKRJwyFXQNLk9BA+Dw4c2NPdVVtMdwDWeWh
CnAawHX29cw6RAJWlzPp6c2LZI0CVQfyZSNAQgPwQalStNxXChwxGWwMD1S7hM66
JkmBYI5/B83eCj4FLQI/b+Ytjb4gGwKkXJBaIo+hMtUtOnv79ZatgDyGQn5oFhB5
GtctCp5CLUOUpedeFrabVIoIWSPEX7ssgoDI7TrHYSFGIJ61tiSbTFPsFcG+stpP
wU2EPkPCOeXqc4RvkvNKldzeTy8IMhAJvIVd/il3/TXxQY33FW4SSdjH54IOmQXS
8OBRN8t5Byui522wqBfrg11e5WSL429SuCCxxFnE3ZAdyQKBKLv7hEV2gaSlyk4O
TXWGROBLyYT9bT4VFYtUHAwd1tfQnOkAc/gFIl0/HTDGLr0jB7oBJ757qwbFOk4x
4Lmim6TzV4ZIfkd0pt6afNOj/045piwc5jji81yPD2Bf19aPePsUri9FVby1Mdm9
+lwgmO7kpnqy3E9ld6vYfu81tr8gQy0Xm5/ZxLKE1KsGGheIAsRjt8qHh0RuJo8S
wCw+QC93ouZYJKhpRXVnxVPktgkNTNb+06FDxQuW2amQxwt1iidqzchxZcSXw7Ih
gO6fIH4XIX8Rj49bMBP+AZYUie4PLUxBvfpYzk8cTdEsOJVYOmYPdQnBTvecmSAE
zZFw0zldEFEUK8DyjM3qYfMbG2Xh/nQ2aYzcUtZaaN8OhiUWPolESlg3Cl/n6uZo
OxxGBv1uqDkP0NPV8cGQb1eI1QE8PKPGur4ImEn8rIr/qhGFwUHNaCD+B2EXgmgg
2LOg2UX8bgtd6xp1Q59yu1jYFfb2ssjLSYOpsIGFNXUf7px7ygGS4KuIhjxbef2S
Xqc1IG1JRLzxxFJi5G+E/mrQBR+NI3TZd360WiKOa2emxpNinxjgk7owlTglOLE6
NMEocBCnPLeT4nctYvlOr599sITK5WvtgsEVx/SpvIqYGD4b/ocJ6WHrVFPVyVUl
vVbEc/cN5or3swq/2uVkhvj/QGQ1TfKc3158N3SkKZPBHQgjXbHE4Iv/2dLWh57L
bs5UmdiZd0m6BQOVN3lppf3vEzWAfqkHASAAQlm0866L0/9neh+ibKPeY/tyB4o0
wUnAGxvgXEGYuXCo7pCjWIDDSrKJHsmTpDO+M3n1JQavW9SWmEWlvzaVCBjjnw4m
SFvQhqdkr11pPP34xXp7t3HCuzRoizHaJCrCGxo+9D3lzKXw08CMB1PT6O1uhmDE
IPor9bTHvWeA5jV/mQQ8YfjawZsMwfchABUlsKm/xLr30hsmPyFDDNGabCH5W/Vu
IynYXvkr0eaO/6EMuNdYaAH40bxXm6GQsLsjpzN15V7bhiOwAaY6GtcgnpDNlHy1
9KM8VuF4vokuVqPU4JFNfZ2nbYxtulpud6BuHJ+KWn7oppcS8P3LPk58nX97Sa1d
hlImZ6y1HpQZL6B99nKAa0bXc/RVjXfi0kxbh2b4peu8OxHXx4Rsky0XkZ90V8cJ
QobLt8SG67ivN+0R2nOO2sjVEF48jg6Vjmhts7RZaDDxE5/5f0sx7SBgOL96o82a
nTRTUTkFUlucImX32THpkOtzqwN7CZo0c0mO7kBXrXvDXOKBP86i0MBXnWrhkQB3
eyANusurpYlgYHHz6kupb6QI1JioLLPY+NLrTbhdMloADYW7crI8hyUd23i7SCg3
Gwqb/iOM3qqKesiSkYzkEd7T4G0xP9wQPAZAk4Xc3MU3mhO8eTfEWnRMNrnEkHY9
H5kYjO2PXL1wr8PuwqyoK1MRU1JaDtfaQQaesFyrPjj3TQ7EK8RtgIP8ofxwxyIb
HBeAZAl776tBfGxSUQyv4UYCNVF7O8LBe0rSBz6YPZQTeZlxLUAmg2491jZoO5it
dfcNcjga5AtJHqMm4libPyWgiz/EolBPUoBvV46lA69EBtei6q7oy1eQRCZ7dbCY
EGDBQtEZxF6Jl1hJLWQvwvvwB58/yGyrL6k8IAAx8QAlWJFrKXsJzqoyRiP2m5Fs
H/M1sVlGbEk27RndRHXkl6rwZnlVlvt/WrK/O1RcP0n/PeYzhpjLbnvwfXYmXdwi
RwTXb+me2x8/eadcPAi0zClVvByXjY/5SZGYrPcENeAU6K8vVp7/pwScqPyDWpvc
1n/mkNETifvzsAB2sfS/FHuTdm1DWFrHewCIx9f6bs2IerjSOHJgJFQVd6EtLp5X
RliIwkoB1fvYtUgcWmKKsF7rhpEUvgEZbgL01J3WY7fBwcWJydVwDbz2e2lyKMVc
1IKdXspzzUDtpk22PyDeTcFpz/ECpZxX2GCjUBq+d8MY4dCrM3ObWSoXOYBEWrip
NBRNsvBWuVg/31l1Zomm0Cbf5fUqRYcXQDIJPCtvdp0CvFCStBImK4/ULx6N345r
mnMMpc/LcL/POmdF9zJEH6Fyp0SzOmkqob7+k3PUYd7UZA9I3tsTpyg1v+arlVdS
qfrwWET5Rm4fxtw0cuV6xT9MWtRu2Woqaa6TQlJd6g6UZ6bv5tZTO362g1qR1VCJ
az5mrb0nBuFg5v5e5hP5jTTLmhq7rGQx2GoWt6tVvTrtAJQ0We00HtOFQXlD6fvN
ZcnFlaHzXOvSfto/K8NPmhKG8DpS+uWLw+XVQgkdaxxlRMml1Fn8fknrBQErdotp
bQy3u7kLo0Da90Bw0ojLbZRSliRAriWe/sm9430W4yknEmQn5ukAXaAj5Z7eYF/x
Et247Uq/3ywclEVzsvAwilIDt5WNupiOJMUZ9puPpuv4sRQ8NTUYNODTB0LJjmg0
AbWTnjgjqXyPcG4ZNLCqT5vtcSwoct/+c9W3Qu8BrZwJ0Dwy0Yj8ljtQgUNzBcIq
SZGUHEZOwSKTdUInOd3Y3O/c7/7BGZ4vK4F0hM7cACdXOKFSMLhMcvgoAl+otMs9
5dMsSESa3SbKO4w23qffNAna3Q7/QCpPITBkBoXeYpjW6mDvHG6bHQ5KaSxo6Ya7
jqD2ldPkv9lPOTNUbv0D3ssYSLOOiUOLw5eiL/4JRfkYM2GZED3bcqTxraG/xNuI
Jt/+WZOtVnoYHNW3T4MD0drb55Zx6sG69eSytz5eJJib9EWRiK3NEkyg2kwHwr+8
8GEE8ONvV3H94ddzSRV8Be5b0jnP5TD5UqERPKYHdtEC5XOUyv7q7TUsmo8lFR2p
QRdHRlxQDKJcrpTjhbJYjIZ0TN8pyCBHSpf9UMYovR6/9p1+gyzcIwukN6FBISV7
In0LliRFTIZYQvpKELF2Bb32IbRERALF97jFMOO9oNNiP6T7fEdvHoUCaMDA2jnP
/N8P2ZFAFK3Vqi68aydhf/hR4UkCHLxODFe5NcSrAxHWy3o+SnQoAShKid9Md52F
AhOUUs8kvoFg4yIbzz7Mx2xH1LKSyFLTQ9rBI4Z05sB0QEvv3VIYIBm/jL61H5+o
GrOdljeKjNU6xVpBmX3U/eIXJrgc66osm5re1TP5GwAMUnYDlwx+zPUs1LYdmJAP
xvg195x2PbB+hjAhk3m0zIxmHVxPSrxfuhogZ4rDGQWKc2YfVMs/+w59WMEXGG7M
Okei+Zw9VdcuOq238HkDcW59YpU1ksB9q5RDppjIkTMkc357myPZPnkVMxHGWk9J
L2UMgYa0NIuydedYQMvtWntQCQ75GDKAR/XvhhRsZj9/KruUROqvz1aN8CV6PUj9
5gzA2L1N1Nb0rb2idOH/Drif8CTBdZqZqmmPjZ4rJrtJSpJUwRqDqaB+aucH68hC
r611YyvRe4q+wzbUeIu1ONzt2JAZONBK67OJfzXEvrY3hyWrKyy2SkG1s5LxE7MB
qmZgHR4DjufDd2tIoNAAgM2FQjiJcVmQbjMcOono2/sVMYuDG8zpa781ZVZJoPoD
6CkSQF567cocdOcX4JbfGcR6OmT7gz5/sIUEeoLtaipafcDesGZIJzTl44oGDExn
Nr+s+JATdMtxnyLvm13CWJPAJWkVBpXbcU/bIO5WWQzDpieKFX6b0ajsdDfYqhIV
cTtNFGAWuEAuZ+G5P+21legKvAXHEOZfBwYA/oxv613aaCIqlK8hsl++pyMvroWe
gqbzHaev0C4wRmZoi5qImCotJ9JGUJDv289FsaRu3CFKOPCmutU3+DOdEtKnp3D8
O0hR3/SpmP4LNSol1tMwcSwyNF6Toheegk57LHZLf/DK4s3OBcJ+iJzwaugszd7U
cAMZGSfa4ol/skUhFM5dh2X0jH2inMiTdKnFXY+PHi/C9NTR0ax1HzDDBnGvM8Yp
4aHeJ2S22mWdXTiEUDk7wmc/FtvVepxupJvBS0xc6AYLZQ7Ols5lJOP+RtONIVLJ
zzBYxunzhpsr9fo1ill0nbWBbKoOEywZZELxSwOYM++sASk36cQE7lMTRVHOxRVd
G86i0gu6SS6KzzxcvyOrNlGikB/CDlCkEB6OTIb8e9c5Eui6jd1frYPgXz1VREVs
2/QaXkUJg/D9nuIKRKDr7hmtL8phWBt/pcl3dYqQWcYxXnWftdCwuIgM9sCS/cek
5Oitlv7mINiCKa8sRuhhphcgjNJvhQeTrc+dmCXf4CHSmrbHbEkDBdqJtTXhJ1qd
dOx1hLzGuoMKg5En91Edk9UDEiP6fdisirfA6vrnzMtBeVHTdRkCYYR/4RGpqflS
FnuoWiVkMGpyJFIgSiD/QndEVx3fWeR8DONHdFdoLc3TNFzY0m52M2yolxx0S7qT
KCbDAyE+JOD81tSwXeU5k2Q9MLo5D8TmP5FN6xO52nCubQ9C8GYDyU+YxJdBGho1
kd/Ytf9la/26UmlV9HtHw3VkYdLxQZw5NrObnL6D5GQPQZa0QDPnVZp1qt420qBG
fEQx3mB4thowXa3oopgm+uBD+jiTbPwpZ64KpFVluvek/KvJPWAhWZf+z7dhQb4n
JVP62aT3fO4y4gbMCWTlT01y6oAxG4b9385b5eQI5/N/qwKogaeyStiGbDbC5w3j
WHG9bTg4HFUapas/PT/qU7QhEKSR8jLguxdL/M91fUJXsaXUyxzI7xm+FhYYH7X2
NNUOCzxZDXgNO3MGEynLPawJoSogaJbRfDbQtsYBms2tN7GuJi0Tq3xMGWNm9/tC
t9WKLEWwFelcyuJ0hI9QyUg2vD6F5dTsI7LxXR+pzagKNZu9NkQfFY1Mol+LDSfC
jXGr5xROooKs47a729YMKnIpe9Km6J3fak044Oww4+kiaE7KWgZpOZT8e3Uu2ly2
st4ScySaH3/6uiHVCl0wtJW310YD49I+XL+6Ul9FMzvlAse1S23hsWnF0hhHzHVe
4U8cvyCclPTraTTI68cJpBEy6XVT6RQD60s+7G9zL3i7r36w8mXuJhhD3vc55rry
PnmLCiu280fZTvTNgeZpypwAxoLfUkyNL9YV1UmDNM+/FgwYPtKftF+Be1E1Cz4H
d0q91B2/6IXSBgO7J2aqH1yPwGwA+Eg+Y4B0pDM9366h7xPzP9C/Qc9v8z9swpfA
RWqlhaGXBmV4uyDpjYerj4nSPV29Zr3IHMRnmSTI7bZYu99Ix31sL2L23UZVtSsy
pZAy+pD2Pmz+3lQqoQnXfdkbfzigXw8PJ9+SYfgxiCfH8znOlwGGyHSc7Yj4GG+7
0XSbPYMrhhN+/FuEBMz4rwqag40r/OIcX3P7jmjlZ2VyyJxEV92s53Ss5ehN2Wde
kp+a4W/lXtypNCa66fGWiyrq9+feLHDXB9TVTSxMSZ+3oFeRp8DRBOpZSd71/UiN
oCD8NS7TrhLV18BaFfxJ8yF5zNWSbpAkQRWiAFrAHF9XvjkMG11HSAxZLxVr7Lsp
g4GFQUE89ZHjT6PcSD7T+yFxljw234MAMR8mr5jzlNQilYP0tsS0XfECAIdqUx/+
EesVuTDZL+FFxNjvg+VuKl18rIbLJBwC1eOZUpnnbWFMeuuyqMtFs5aLOcErxWE4
n4KI3vWmJbiyEUMrod997l5L8Tmri3Ve2bcEE8GPu2Nxbb4r/I9sa7+PU9o8dw+S
oiFXWGQwSeiQEbket+yiFYmsTQqfcH5SAH6loUBt5iMRC8ZfCqZnJ2lJon27dez/
3Z3lUfCrKuA9xQ+6aoJbtxx37NfnqXbO1ESxiwHKSoVES2IQUd6IM0eMDHXSn4Iu
HLBUoMBJ8AvRqFFAomqKgKbNJ3BxihHqvEpPCMlUUdWt5fbCNbVM6+VqYmNVlwMI
hRCrFz91nnGZps0chWl/DtoW3DPwvVy8Dsl5d+A31Fje970k6zfeVaFJ5vdY1S7M
3aENn39OHDtQOZMpgS6gxNnSpX1dr43cd+RXTK+a6WyZUCyUivtU/HDN68E7kD3m
bhdrvZUirPG39jt8tCEerh62WEFEp4aZ615WzrfY5Iv4dTwAwBYZJTch2uD6MobX
IErqpgVeJeN8rnMy1ItgSJIB0gvyxcB7MxVP1SKsaq6AfLJZQzhCpC/F7rMUC2qg
/mSC0ePHoURO4h+y1/6v+WkmrajeVggSlHWNWJOTEngXU17qfNfbzEP5/G0AXcXy
cjWQupE/tw3I1nMzYxkTkcim23tFLUs94X9C7+EoREBa/WTNT408DqjRQJ1/gBSr
tywTZH8RgJbLHRttCsXP+V22ktrsR8Ho9FFg0QQ0cHteVvqBUkJ5jNPgbt+HAWnj
VQzjBx1p+iFYLLC8/EJKb15IkODp8wBqxiUryUKKnI/lWpB/8KskCUrLwVwGShgH
z1b2s3IDEcZbNvNGyTPn6rR6gtQ9VSsVnDcKR+BTrwbg4zSt4E49xmvRsFYfnFhg
55CDr4BtQh+oRVH4KnXmMeuco77FpCwQNmiZHQj4VT/VkNsUsmUWr5sz7uH7PDhS
5wMedj1lCWHV3JS7hHQQLuEIfH8jnT638akfgIlkwDOFrDFQIr/BUPgNI05WvYfR
UWWYdrnF/Wy3LVYyVFmx3o1tQgV2MwNfEdodlQWVef8IwN4JYd/qYN7jPqVu0v/S
MMrlIU0SKgr2l4tvdeVyliUJrnwUFwCxWGFZtAz4nRuVfgEzd9N1K6pss4qHxMTs
t1XRWKCbuXObCwoQB3BOm/bZ8bOWL5Hm6mgQsVQhqwNGD+km3OeW7ppdHMcZZWr/
RvJGsu+qlLp37SR6Jz8va8OaNE3aBlcA8ii1GMVJMaL6StmIDKDd4UUDKaMBLzLF
2KB8c68tDukQ2saXSFbvT8KddYzNwpGDrBsgyAY/Vayn5Fueqij5esB8p//OVsKM
OSIPbEwqWAUe1O/o50m/3yJJSYU925ICBT7KnzUEQuiKlL9tKE4tDYRNFqD52DVc
mR3LMlvoA+DCe1sEPKXf2KH/+T2EDeAoc19PkP2+0iHt7WKQVrhdCTsgvCgjG/mr
IqrrNh7pj74KgMJB0HgiVrzUCJ9nwyYo6npKUugnnsVHQiT6TB//S0+BFThQUsh8
WKPrEb9zCXDpMXq2Zq4BZf5+Gn1YulXMguaZFjr2V1nsO3oO3d2YPfK4F5lqy1+w
LCxU70Buf/sJ6g41T+u2lyZtwOtXlUNyZqLFpxc1nsBu6m/wCxUTJoyYrMWVCULF
P2A98qm/gkrHextrWaZWz5zhot5daJpyEIiu9SKCGiOwyvsWSceel8Tkaqopei66
863r0Esc9+MtR5s/HrqdW/l6aCLdjhgpkhDTfXIcdqAAwPiDahQiSWwCts7zPsqK
KYDlQZ01NaUnI9397gYz/lfYZ4mspJgtZspKWJEVHJLwLhdTnjfImlaEuVaWYFvt
WlthGsjVUJUm0a977cB6TnzD+lsU4Z9AoLeL4L/pt6k5MGmDNrSlUFD7RmCMvQjV
s/vwr8WYDsjFH4fG0ZusSRTTaA1xtJmCkj+e/piwteNdV+KvBl5DBb4Cb7xGet5s
XGp7QExhJ0CgIvljL3wLto1pC8d+XfmAYNd4Z0XhmS6DbSw1KDLRyv5m6lRvMEY+
iNf7iZU6ZztepH4kd5cHxdzzRM8x9Qyko/3sKA6T7S7Xl2/tpcqN8ggi+CwQpdaE
mw3aZWrXRQgNqftWKTx+mQJzXYevV8Et6zG5AqHIRNQXNnPM34O/LewT3hCTKVi/
eBaXzX0W87TCFBmsTxhpnegtCtwcDZEYCHAJuR7l+Cr1u3RdCK6qU9LzTwUoq2px
grCv0XZLLDjsdDNyJnjKWeLc/xSbXg1GjSqeS7bizST49A2FaEaBZGFA0PV9Fm9E
06MpoP3TpmFMAoOwlcJGTntrOAccVAHG4gy74wa7Mb9+0e3MR3SuYZo3W7GsinbN
/lUSbVPg86GvqL9Km2PBIOHhUP8vp8lt41oFink5CrFyy3M0UVRkDgH3HDyh+eL5
D4Gd6T0PFbPEM62vMktTMe2EddlGMwi7ESpOdobVbcFV1R5rbwSIZYvokh7JvLLB
aKcFZIWvNpkEZlq2eXVOJ4eKoSGAaLQZlYq0Sxwgt/IQDK0JLvFXL5D92E9A7g5N
kF4wVgwh+ql6p+W7gLQUpTTUIeEWK0Dpr4YmzEz1OU5cUdq050IulmZgnoIUUm60
jKuKJFyqvqAOBTGb6TRv1G1vFw7ox3UE91nmoI1Oj6xWUWwu7wbQ88zpeaIdBUFV
yB2VO+oK3cI+fv/LqPo3hA/tp0L6uI6cZM1PJsDohNrIMnShGTc3hNiK6bJkcrax
agiw46ccKx6vzHBijtKnVejKHa297CvD4mGpGynyYM5BsOEeV+/3P/uphuYow7HA
OH+nD36bJyNI2sUXQ/dzcjovdlvAhpZk13TbNUQ1mFrmO2/wrPXnpLrmHMYDNDge
N442h5mzkCt0G7vIM2jlEG994gsFCeQS4I6Hi1jivdcotn2hFNUFP+Qbc6XVtpY2
8oeY7lSqwQBKcuIyBfDjfFzWGlpFwFm59R4crrkrHA5vz5nC/si0DM6dCFQiNF89
Zbb+C0GPIjNlL0Wx4EjcWvhjMVqlIB1aU3fUSUwONVHJvoDI99btcUYwFoPT7SZq
GbFnp7HjK/SbbYUugLQGJlj0NgF3ZvxarnQe5j+23jt2YsGzUibGiTuE+S4Y5Tpm
q4Jw4/x8/5B/o217RUM4ZQwDMbU+5o+iwHu+rQ9UZGGYiU2O77GLBvErS1vpROEX
7uCT+uZl4qhevUBiPeRwtYW8up6+LLZuqD16Vg/PutdapBdrUN75ii2nI6LbQKni
V+xyT3NVl2jYDzm29+SgiersO9thYiE1RyT6T5qvRSkv/NwxJJqLomZr86423btD
aeHBHq7ey0QVVluPhgP2KH1z4E9fAuolRInqxP4c9WaNC8OKWSa8hYWEIvHvKHzv
oLU3NSumtn7BD3uXnCwCDo/w7s9QTAWK5R0+mlFuVgDvX3M9wMHSGXlWNzzXckdr
`protect end_protected
