-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
hkQW+COSm86x9Vva7vZLMYXmNaCmkegqiuACyx6ynMrQh6Z6qKQjLK/oSy6XgYHF
Z18wVJrOegjbcvrtYiI9AqH00bcVshbthFuAqy+adH20LoD7MKhXiYgNT/fMa+m4
zddjPaYuX1HbAnoHyw+mSYdWJqMRE1go4e126JAp6YA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 7808)
`protect data_block
48wvaU2wEHWVrFb3GScW0MA7nNXkWN3tmhDFTmIjVjw7frzkDNcMw5I6U3N6yb3d
4+/F7xJiD15t6iVmxj2Rma8gmrR8cz/FoF8e9LYrTH1wguipwtpRyOOSqaYFgYU7
d+PNhkBtbg2BbI3NHi0VoH3227qm+dQyWmp3ADYEOo7AeymwN3Vkwwfwr8XfINQV
YEQxuhnUVoKCiF8VpY2xlADf3L+C47qJ1P4y/dYfQL9fwGUPXtoOzzO2KKhdKlm4
BJAA4/e2Q1a5TmHJLXjFMilGsXmufHSnd2u5QOrEBZdD7lF85BCf0l3vELEWfkvJ
vUDZ2KOrFJf+zIMygt5zs9SxUKzqC5G4ZL2ptZ7NUMAH6cswzprTSUwurIMGqjb+
GrrNiV1JIUsa8oUtkqy5IVVMywozHeLYqeMM6u0pr5VerDKT+VlVJDY51Aqx8yM/
8xf4ekCqNm0+oRLZO2VvL9mAf7+oNJlkjCyV27vfL83gGvGWiLvAJXoIhj9mUyLs
/8YUKR8es9D5KxxlFvAGq0yPybeHEEO6xMCc3dPC2xbQHkVfKFGzQ32/gZECkBPl
/s49GEUJ5qlcnl50yRQ+ZYs2yvI2X/ziZExrj2BE7pA2Bi7eWkT96GZ7jRD/S3n3
Q7HJznmEUVrn+UI1t295m245lGJI+IC/FPZyae7bSAzbaqGQ9i0Vsx6DdrQ7rTZD
o1DNN5eYTlEinbYXYnOxLfJtn++PWoqRMIAN0kIagrCA6VAM5KgtcuL5fLXGeLXE
t7Thc/2uCq374e/0J4tNgmf9ds7qebXZ5xmrMNkcpFz6viYNUhTHPyWUEUPQmwxy
vx458NMq6iRNKsG8kHjnVmdIVS7zaX3QdnBZ4XHsn54HbtTQIYxNfpSKNo/5zdDU
7+09qnrNbg7kWDqfmJDcQ5uwtPZ0k1BYRg2s9WNYiVQ4VBiuOZbtoHcbU00yyjdg
B248vDY1OL3ArMx5MrVbXW0kUG9PBHnnMKAklMCLaN6BS21SVY46+bsygjFNvs7j
JG3A25rMjNkB0+Qi9km6irByplTohBsm/enRxOVE0fIJ/agDH9vvTZd9JgLwJR+Q
yBAbBuFC0UjnVph1Grv94rqOkkOj4A+AJqPeYrJBZ6JWhyp9NhHyCerZTwRsN4N5
zizVSmuDFMMXl1KGaTsb6yGNyesPOEjU7w29uUAjTIRLpQzBIIfQh3o8XIO6ZSdf
b47sasGXzatP0Ex3yE74uSa1ga6SQc5VUb+Ngj10qLogGH5x0iL5KAT6ITsz1Mr0
7+e858ZL0NCYOXyzndR6LgSnbysl8oSgdJkXsJhxnFW2JHXjqGmFoGAEEO6jB/Vw
TJKYCxeUMS0VdCiXN7j9foM8/dhs93mG6Yw0/RIbqOkvrdC6hmFntwk8qbKN6TtR
wz6ZRbKfaeRXupVp2vMJd6oeBs6Nh0KEioVeCvaRTB+yELRilglx/WXougwXtoXP
+m0tUcKKCICOLPyfRtthsXLgkoxKSKTeohb9XSi96kCpj+RRjohJog0DWo7DeBkx
CmMXwb41o25sloHrrZ951+7b8Kl2wCtNlB/9c/Wo3U5d1LI5Vzley7GJmFDfmJ+G
nqJfCya6Qxz3+xfvihwQ7yZxmhrNmUnA7jdlrVqhgR8JfRI7ejhsR7tROWUuxvoU
lJqOL5WuasWKAWxqeHoRy+3wLcKJgzSL+T+jFFc6EHWlK7e71/BtiHOwOoEWDUkW
X/Dy3BZMfBFCnaUGdLzSW3hETNBwlwM7RJLNZHNEmtgkBYBaM3Vw4lK75OOMGhol
AKV+EzzhRwD6XkfKZ1DU3l8lT2EFIdIuCXJTX4ClhqqFiQ+qM12dC/ZDp8mKzWqG
q2TxRRO74RJM8v0BpIa1gml6wef0DLTKtCvy6KNYUW+6wy4qavGgOOckNxAPZbfB
EsilyR+dbyE702JR/3outui83oHbdkYyET7yRYuxiYbUbu+Qt5HUnCXgZrtiHIjG
fNDqnhIOPiqXaji4JpodSOTAwXdfJB/ebZeR0t70u1pc9MSbucL014exIjMzz/rD
vVeS59m7Du7pTJIccPWT0EbyGc6BwlFMKMbsuM6A2Nzfp7D/qrhdw7TYdQj6i2pt
MmZVC4P0n9QcxjLshGdUYNnvyg1XjjH0uvaWImcILw+4XyvT2dE3iESVAi2KSoht
fRv4cwqb5emmnUlUgM2KeXp7et/3gpxyP4ITW7F0lZKVAxwpmAsHJN0sIwfc9mht
3Z+Rwa+ESqZ1ghtC6aUGpQofJ2FMWzvhD69aFgw2guLNqltIkwPm11b1LkVwMz9x
nEPM2sjuiEvEeiyy0UPC4A9IX57nYSUCM9Wls/AxRAihWj9L/AhidYou6fZr9WN+
ku5mOFOF4OMYZ4hMBt1kfADFMtd9/iKmM8MCHZAor+asFHQZ3v+sB/i84FOD4veI
2DoyaUSMaUoHWY3Briten0ABkSWtGlEABZTx5WpoqgEA5TNhxUUz8nlCRzSQYAs7
TUJ9PX7hTIwsoyS3gVq7I7lGTiMHgtyTvmGEexegjkzmfqRhUi+qg5lVGY0UR4k+
Z8QSMn/uDKmfmFEjr8ifDSaJCE/SgIJ9B3Do+98a6RoPR8UVK+AqgAQ2O9S2v+/n
CANifAxxF1XibA0jdDBGDP7Or8uwCx6Gimnru/Ay12Ec0dkEoc4RPprYeoyJg/bg
hvTv4DbzIGbd48PaqNVcDb5L6VJ/VmmoK0GslJ5FMQV1cJR2FxXc/j6851Ucc7pr
vOYgu9D3IF9v0N30vZZrGAKE044FAwaLOHX3/+dZvJSEBaJ/5Z6uPLOez4omOtVT
gkJMJTtBukUonCwjHcIeM2jWjzp3DRdzB9xu5AJoW9evTwgIXWlUWXMCVHlQtZzZ
VnEOnlW2MIsf5zV2o3Mm5fAqeqOClOoQ6dunuL3f3ONDXyUticgX/8IVKttHfQ3H
WBB1G9pQzyzW3Q/nJEQeHb1JPa0J2/q55p2I+bS51U5ABPr/4Q8Kn7xFwum1KCFf
53gCIzu5BTVgbpNIZol/+Iz9Xt3e/Qd4NKWloRMykrV+M4JBBhENq9udPECFFhHv
me2QL6gphEA6p4mTQjb3dxQClSEgMfkZk6dEeVFsrf9qCF3nEuku4PxZR8KzgkNa
x+CCYzqw4ySpNdqd7pckM1LrFqnt9azjdOSYY+Eau1ldBEZ3JOxJsafhK0Tzxa21
S6K80rNQfmnxjcfEnxlMfCYh22z17hTPKYonVqb1I/aEkOgaeOZfPlX+IBtwBlNf
bn/6PxZ7ppXrG38kL/8BhWwoMxZruGprDJcG2NoB3vcfZ7/vWqTKIg+gstbxODhI
iV5fgzfUK0Gdy+6eN0tLy2pWPG8HDlcExDob39usrR1e/TH/50DGAQfXKPJtOlbu
eym+jq9uy3NfsqDqO2edSwN6o4wikMfg9wcYr/AtLpoLAJSK1gr69gTQd7NBgAu8
pg3yoJzcC+HB6exsyluDeMrydNJmA2lfP0ewi/yO3LMNSpiwwiqO9erFHKgcHYnr
sSNrptZykSl+ahYNdLPyAcqHEJndrmc4H08szpGALxQ7HMzuPhwOMyvgF7duvgX0
O39Idab0Ba2oQCs662cZtEjGnm+81ft2p6gnFZl3Ao48jmnUG6FuDc+wgL12gYkf
YzII+iFKKwK2h4PIBEArG+Qs+utn2RRl20QutHosBby242KUxippjh64KvgkxLre
5wnitDwM3zd1/bIO+01fR5S9g18JH2b7utYEqpej6AzoCNkXH/8oYpiz1VQvkKMr
/t5c3ySRDnOhcsPUQ+jIwwh4vic5jsJEKm4aEicic0iwrQ85pBfij7zkSTn+27RO
IoAqQoxTBXpGTSkHF8Cz2Nh1/7Kk4In5RfmU/7MsdNn2a/q79IVh2q/LW8G7VBjk
KpMVrrd9QxAFAg9G11xj2NQPgp/e0/5RX9GU797AODqKoKIxUDQlJSSDtICnhNtp
zXUnOpr0QpmC0WPRVjZW/NxraN4TXs7Z5DOYu8k64LnGarpSgoZmNg8WilOpqJQk
ZzZwY6bEiW/QA4erpN0ywOL8CpH9gadX0GmQ0+WdVMJTdiSu5WiXgrXmtmB32sz3
c5kHNG3GxQTlRzQjHI9Ih+5GK62NRqN0bz/eeDhANHkcptOZHxLUuapeiXDWxfLT
5+3ASxXLyIJLM6NMyDqwM9kfztkRsHlu7nISWbjwg1SFyauLtN8kP9VhtjC70hw1
dfQUVD+AptdAG7O1VgPJoa0jB/A2b4GfV8pzUAEHwy8CMWkoFKK2055s5thoAFg1
/OuM0QIQAjucmoT5eoMmsWdB712QvWdgLt5rCXnnb+tJzonjH8fUTU1mTF5iJnqW
ZOZGcpbiQt23Flx3/PCoEn2G1qtngu/fd1FDf+onKFtaIJlGdAfdfZ+SC4yE1VAA
GhrPy7uzp4Lp4DPF3e6ztnnafkVGm0f6C/CnEGTKf4h6yHAnues8HNRe7wv09c6S
Qa4+B80PjwWwBU2ABPHyplVh9wuG/oWHU4ZxBIziq/8JwEFU0nRc/sr9LTJg6iSQ
4mYMAkbpcosh0lwWpsfGAPS3Gyd7i/aSd/9QaeKvt6gYAdffYeyzFd51cEMuaQ3o
9bwJQQ5CrL369E4wznHMMr+A5bppvFTAx7QqSBRvb8I3O19el8RrFuz9b+8x7vmA
4U1uJj7ka1FPJ1GWsZrtowAs5xyB9LCW6mQDWljX4iBOcJAoZMG4L4GG7xvSTLZw
yG+8DkpjC+jIBCJ2uBa5mBmUWiEXku5eW/9P5OLEy5m6Y3ATTY8KogAjZx/BoNgv
wN4mhF7k1x1ZjB9IoPkCeqZ31q1v3IQdP2ROHQUaTEgGmIshq+HhvtT0CWFa4tu2
BEfHIp5/C443W0Bf5WzRv/3COlhXpkgaI6i735m5F56vO/PfGd6zfxsbJY6fB7Ld
023nTlCqjxggRbpSFkj5uh9k4F6MTGoBEaGnulIs36U6Pcy/HkyiPEx2wpvRzd0s
QDTAJzTlbg9ZfxyHZYayVyYiRLDGXOJWf1gaVWVqJ3TBekAMpOn+JmmlbN5CQT5b
V74LObO3pIoK3+W6ZpSc9Qlg9IEaOC6WXyfW9pixf89PCk4hN2k0mgQTg38Rxewd
+ykwCkuAGIDk9soGt5hqeZCEeUe77U7vmH8d3anEE2esRsqZiQC//Fh35yCTLgZZ
A7TMCyNRSnksO3tD/eHrxwjATxsDkMdCLl6qLw6vUU3TEG81Je5uQswpDtMCb2gN
PeYDBoTNHF0Q5gRTC8zcEHKd00yonPSBrjfEwVHtfeB4KtQArdLFxQlrp+bBOrEe
c0hfahoAs0WFCFTHx4B4ytcCKDJpUwFwddU7UqoJ6jYQ/wTIeyPWsfxuf57+ZGNY
nzJXe4ho+Mll9ORjuOG5fuK1IOQPZ+8P5pQMA66R2qWbBSScbCbmAQZt3PAewy/B
hQR+wD52ATECBRRfu14MeVphKQXARbmCzDb342/snH5OMzXrJtjLaiAu3Jqliib0
+mGZfS7Cr4d2/zvxQxztpsoz+q5dkxayKqdEwFVQWck6LRYRGfE3wAQhO3JtsHlu
PAl3Em2573ffCkN/Lx4RFkaQO6qCGfMRvY3sUno289zmE9OMQm6I1R20xhHUt4Pj
kJ7Y6AsXPq8jAhpAYRHMVCJLG1Nn4thI6kUKiYHIaP36M0zyTSDLYA9xxTpODvUg
mJ0aJ5N2qhX7f48w0MAOHakyE/rki7Zjc3fVTfsF3TFiBVI3CI1l5Fc2TbU9scJ/
Xz7kBgSxajL2WI6y9fbZR6F5ShHk6Q+RmXJeXjXe/L16eyOgNBK4bOu32Tascoel
Zh2CJeT3wKfkNcm1HewHcrLxIqJZUHDtST86XTtM2qosMq/V7kK8dpIsHr0SJjKE
fjJFrObIoYY0YHR8meZ+dCIngKXNl9Qrxt1bEKwzh9P4cn2esENOGGDY5GGA0FTF
yvi7sjXZC3sjzlAXUgI7lB7oZC/BPraQYRYZeDDSeItz+qzKf1VEzfWiiPDN68/h
JBLsAP6RtSk59AdMy1fK/rv9zM8/5ZPOHZKYUWsGeXC+y0mYO9HpKp37LgHTTbea
bBbKhYwLM6UrsDHpaC7T2D+ptxj19uJqQfa8CS+FcFjpKaEqBXPEcozYQrNx5Sw3
YB7oNnjaZSuxOh85npWbSuS43INlk3ylppAbl+25KUrKoot+9kNYcNbDemHANESL
HZC0mSAbZWWXLW3TWTz+0t9CXpi3jKTOcpQLKtBQzJD5XX5AvZrsl5ev3H47imFy
cYIBn2wUAubIdFcMWqZEU+fvdjjgD4ZfEEmuOu9XR713D3voK3zA7Rg1VfuI1l4m
AxdS9RGkxvn33p/eebOzfH4p1J0Tbz4hbMqo+wlgbcRicP/ZzOCbT9ZVr8zE08Ss
CbQezp14PRqpVcX67NizCbW7WiVdYmMxN3rE5m/KgotEE0MP4UR/mT4GsjfOHmSs
Cjj6BzdqbjqfIiF7KmVd+HQiEMbO4mfEGoseIMPUDXGLiUvbOHWfI3b605A+SomZ
QohXllQ2P6SvovXKB23TXe2ts52FftStRnod/whZh3zcbuzKZif9fFWIeJXLxyHc
tRKiL8WAw5h++ZDqDYCN8EltGuOJ/hUSH/qYdgN9WHhlWzglSY9RtY6cWFjpjUUH
beooXAVW+e8UPr8MUTojmdwwU+UXYiO8qsFZQHpjd9YHByZgr9hVYZ5HopiVh3WF
nI4U08Yoq/A9xwAzubHoZt6WS6H0VNKb1BrKCCiI4dg5aW0faTBJ2wB+skGgv0hz
lTIdimceb71DnRsxSY+Mjt2+A43eECkvUspNXb1bVyew0BrfGlR2TNIvIxJn5JJo
v0fcy590YdsBqX8Q6SNjxkcwYHOqnk3eYmW6ygjaMzgDrsQqdDmTbQWWucqR2/+o
QSTj5I+hybvJnB55pbNCEahbrxOyY2HU2KDFoKxNHpJszkfZwFUwLEZKODvnnx1z
rUblVDDYHP019QtOnXM3ZCVR18IJ6VoGGXEups8WshEmlp2ZSS7Ybel3K0TVd5mk
xB1IpqBwJTIYgcWWPyeS9HKFRickjdjCb9ncjhb71iHap1/N+dozScQh/hb02RO6
rHMfwKX/9CL6WJ0rnBHzMpz9B/LjYgie8VmwrVDY+oIZFJuHqVE9BgoVRSaqveO4
iGwLLdHSt2gmuzWDxUyh08h22WSWYanpfQOxorJqQij5gGcwCJKoPtFUBh19c0cB
QeKoMsBsimoCZyL0R+pV9mN6ZkZEarK981WihV+R+z20hJIFavLU4aWksGPt07Yc
oaqvM3PlSrfbWmqbm5+1Frdy03CXZ7BZn4FRlscrWoBZ0ZiSimwtZj7MYW4IkzqV
hWAUJvGQ2grPF49e3fNMlUHfNHxh3WLA/VCfZeEQ8tJrDjNgYGPTuonLF+IOI5R3
nBKnG5zB8JaJCWH3o5qzHKEKgCy0qeYSLml1BtUTQHHIzBktAm5orEq5zAyIm5MR
LOENW9l9ozcUlPLGPz38+dfXeByFiPFaptiJvs6EkB1dfLCDXTMJ2HECvUDsk/sR
HAYiisA/066RQc5B59S077s1wK2XVCxeBw/xM3RyTcXCj6j7ENEnILHIiUkTOHm6
884AQG7SDHETDwr6qamnlBc+nlzKIz7dgtbzE1uXuHnqd8Vb7GMliNRlDQy0PVzX
ZdxTCTOGClmKek5BvL+LTYm04RV9GAIviEj0ZxuQr50hSxnmWM60ere9T1J+6f+T
rumAgm/VVDG5bldGt8DQeDJAeO3t+OK3IEa2jVDLRsDQi1Jczc9JvdZU3OyOwZ6R
e7sgBBOBI85yPjwo27tsuQdQYPdDEGCSykIPE/fJLG3b/7DQkbWkOif697EX6xGK
slP408IgqIZRHGR3Ezr6CUIpbxk2HP1pBoWSVxMw3rwF6jcpk6N3zj308ERnvPKF
B6EhRpsfv6ERdRKfEcTm0n9XZ0tFaNr0uYrxU8ooj5lQq4ZpzY00Gsi7ozqlZCcr
ql7MYEhEogk+wJKFQuI17NAmTE+lFyxWSqtumG45jej0TZcn36B0MP16lvNslFES
DMP4wj+o2LfjYRkJ1D+P1pOkd6U/lFIQrr5TpptBITdLaDRqER8yIo11aX3zrtoU
qGRy6Fxgq2PC1T1fQletd6ruAitlOYBzco1rE/N7/IpKfvEhkJS8ySf/9TBpZIOd
+kyHrNc5K2bEmaDHifpbE+YRYzqTN45L24FFNbBT2wnbRd+Wmb6+9wP3kmTiqDg7
16nVm7kVCwZf09SWhqlZeTWSndp5aR9CcDh9KMOZNxiblsO4acHZc7nt0z7mLwAB
OB1m3ReuTZJgVuC+DA04cSeIgK1tBs+5C/c4I/dgnWMPbS++PrfvOzMdloVTe1B2
cPQPT2WIpDG4oBj8hu4JC8m8sPSmu4AJlyjvoThOgbzzDJUFQUahNGOdx3FBp1LB
7z/e4qn1RabTX/15ymrGvKaFMBmDS/B/02dnay1jYi4+9W2WqJHMn/y67zDCYhbc
jrHFXZ1g9xkjXzr9MpuwZ6nuJY3P+B6gdUdKNkRf496Zfvy8sEKaiUkn3QcLlWVa
C1t0HuH1KsSn6geIPyNKBsQDSitLFiDHscMj1WjyCjzeL3z8kPIZNPrqb74ePU/z
yOdp29InPTagbbdCPxfmLMKc7zL0+q/QW2eQyv5wtxqTvzDyhbRTl+zoay56kyt4
AwjKrl/eEEEMA/xEe6ybL31NNeKA/V2qAMJ/YYmGiSnHHWTeJU4arGI2VdgyTPer
pYhDeUoIuh9QpdZX1keF3mXaFpA4tcab1hDseFT3bKvFQziI/UCWM29PU2oqB6fB
MY63/2e0umvyf+31JNBMWZO2tgVS/CxX7XC6s+Pj2wPewYuJhqMngtGmLYZiYSGh
PIqFOHYVS5GNGqubtlxJ5Vbm6zk6R4S9z/mBS/SrSaJMbj3El6yvjJ+kD41Xbw8g
w16KFGcM18DoBddiQ6KJtyrpwbOxWXe0WfAuGQGHMtIvRT3kPCalCPTuh8DmvADw
BahXK7hmWQy5hCq8yCepbYZQz0XfPEoeSYhcK6Eg9ju184P1C0FZL1wZxQ3UTobd
yknGhE8I3Nn4LYOl9YrfdETVxwCqosiW4sQsuE+qXOibRher992jjD8WjtvDJeGv
arZUPpZx/AS/HNOGWvGSWHzfJXQTjBaxni0A3p+xQHWebvuIoOVS491MHU2aSOXq
scpDJH8P3AKrUarzHWShmnnJXHV2NuZJAMLGuUF81WMi2gZR87yM2PivxsujzjVS
woCwZgzDkIlFpSmmyoq4j+AbCEUrz2zYlJpOQ/zIL3vacCeT/L74LUhfLAxC9ZsB
5nlwxWLApigD8BsrVXtUVQdoETorWVwQsSX+FQUwzOvTxOS3+7zIsec8LoH/l22B
d7Udr0Ef8UR9yr5UTp+JKKbpEGu7iK3pd3faUn1f3573gKQI6B/IorCjiVUMD+Lx
DwHbWf+/EnsgkW0uJOoclbhcSqdChxqgGEnZZDpKAEQNHCSEymIi9yq40cxNmehF
AHdlCASBgrWZ5LVMUmrZsjYUbOloc3IHNj0SxuuFthz1AHR/KWyuAAhOTWXM//rX
H7hKUFzZMT11sOT4FeyCqXwOsiPyoqRUvvXvqFn57qLWjEHKrr0YK8J+10Z1qyvS
osuUyOQWNwXywFdiueYnprqoCu4wJOuFM1twvdjZBuVXJGr50VIfimcRFdEZr3P3
7ln4Fx4yD01EXtpQsOsKm1pMGveWrZUNXsvvIgMcDkVSHdbwV+uCbu3rjcc92jKp
6YCcBnGb8ReQ3JCk1/l/DfvjACocxvULzHqKiI/2CaRxQ/mQcAZ/tCZpEAB0wCvV
r9zotHwggM8tyWC2DJcMUyKN4jt4mZLSiTCRbNwbdbGBnDDyaFfmmyX8vf7bfoOf
wXN+uHYoyx0m+Mv7otqVA41QXIPetjlKbVP//UJ0nf85ZwYNsTPZfC3p16CCBtl1
QI/jjJH6YpOc3zzyqy4opOf8nQGwHxX9GgG3ZTddrMuVc1SwxuZLR8myT6WQsqy5
mYDgn1Rn+NC3HKS1Uorb+oYhuPcPYbnMfj4s7gpAg/+QgBqm2C0FFj5JZNsiEc9M
ZUzvEeeSNtnQ+4PHTPWK1uQY3+/cdXbBROTEOuZdKZi2aXFe2zmCYZX0SWfjRbzq
cl2XQ4Hr8K8vgFBOUAINaQagG244ZDWSydtmvAOzo9RxO9BI4ozv+qrG4Fo33unQ
cUD9tSLH9eoHid7T7BG+7HDFn/QqjCS0+Io8wKU8f5gECLhrJlhH7N9+JxG6UsY/
dsWlRl8+VHFhCGkNXfXztAuNiu4fXn+bi2Xd6ZOTcplPZEouz2ZaUYaJhRnBqEad
S2f4gXWLzXyoIaQKvwBATaWUbe3htVCIgaW9Yy92sFs=
`protect end_protected
