// bform.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module bform (
		input  wire       areset, // areset.reset
		input  wire       clk,    //    clk.clk
		output wire [7:0] q,      //      q.q
		output wire [7:0] r,      //      r.r
		input  wire [6:0] x,      //      x.x
		input  wire [6:0] y       //      y.y
	);

	bform_CORDIC_0 cordic_0 (
		.clk    (clk),    //    clk.clk
		.areset (areset), // areset.reset
		.x      (x),      //      x.x
		.y      (y),      //      y.y
		.q      (q),      //      q.q
		.r      (r)       //      r.r
	);

endmodule
