// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
HCd2kM1f38NqBbvCK4qSiaxLCy/CfFbDr+ZsSckOsgpApcqCboeG0yxgpTxxl9dV/Osu1QsmLgsY
Mbksjx33W86aaO0s6BzIPyd51jRhnJqHom8Wv5L73tmCcKcTTRQ4oeJ4BfEZHGgtiLJk21sTvfT6
sLtZ3n1vb5kDCfXrOfuWjY7k3WlJT4cxDH9LFo6nzkC70Ly57imRgdeEUg4xwQaH9m9689lUB4/a
IGnrE8Aip7oLu6XIGJjEKLoSHXJIPyfK3eQx567fHDrwky9Wf1s4Gi0HYHhBMzQhDGpu3M3MoG2t
DMWyqc6+OjTIBUIITf6pBAnnQ975s/bXqUJ74A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 20544)
QbSFObCyU7brXzXfUw3Kq7S0gmcydvFj1vw8HmwHMJLOJ0J7zoSZmemxL5IwlFM3ZFX1IG50Nqoo
ubsP7hD7vzJi0G8db9miN+EG1VgyvBs96mOmFL/P2JyhPYT80dyOEt2jr3DXONeNrmYNye/2qUcL
JdiPiZ/EWhZhTNoMu0nmnfXaRP1oql+Y+66QjawkDXsaAzhvDfQYv5DKVtAz8Iq9dOat/GiZoHbd
EARuaRCGgDdgC7s85cncZLsyXWNVln9cIxWSgQH327lpShRUEZj+syAhAG8nUujQ3dzYUIwkMWOe
7lBXqDppj6whiwIIxeEuwakObmyCOVwmPhpwb8Qr4MLYSqKQX0D91LEweGEN0iK9XkWglk9NX20g
Sv+bkbmfeGJ4r9heDcfJlFpBcvDVXX+fwYZ+LzqibGQeOzJfpk66/54G4X7l3eDRyDHFnZIEjkUw
WEU2eaTALUtYZkvr0eMe+mrz6qqMenwSRqbycLuD7wYQ0v7wM2CS1b3qMY/H1n7h/S2SfTO0VIvZ
+7k68VsqnF1TWhwgDXTFBEMANEuX8X/POf4FF7+xzFhmxYGHbDLf+yy5KOW4lAnsR7Ucvjr4/Edp
hGTVE8oskK27sAic3RCpxrbY6cWJvsAUP5Ah5tdNQ2juzdPePSOnP2IlYizr0GdTlS0ki6NrOPLK
5YgZTQfnwazJQ5a0w2I2btemZ7KXDHu64RXrN2PJS+6Desk4jAo70s4XeLzHXy3IPblcD+G3ZcoX
v6puq5VYlw4F0irht5w4vOVU0PmYPE72648Z1dAWkOaykAuapGlGNja+2LOw0AvCwSDHxlUneB4o
KYd0hissjysDF+acf2wHOu7uaIzjJgZw0b2giSoAC0k+ztKtVwHGICFr+x+S9wZhuTzkeuhbQXNq
zMD1YyV3OZ2ga1crVijb2xpHp7ic0UaT2gsZvkiOwhrzfV1Go4Xx5dAFacQd888qZyenfxGmVa6V
alqAOtrb1/lgE1hsf5Y/rwkVnCLsXbaz62OoD0v72+MWhIZdeX7vVwacrs2hQww+eptxrX4Q38BY
Y9biz0QiPLpcW+HL1Sn/MBjEXeXMpJkCWNOl9M8/rbZzHUckFZ7pvHVU8qKNWatoPuVAd4OGkctw
kVma2hCu2bDUqxW8IQjALCUhi4pT+8Mrd7fT05BrjKJZRn4jiA+aZvT5L3eKq6xQ6SUbZWCCmHVn
SGEVkAC1jY7El/bcXh4TXGt37Lqb0z60M7KjAXKh7c+QwzPbkmigkGbOFcMuNfImSvYN8b3BxYlL
h2sqiIIRD82D39K2047iRN9ym/St3Tb3xWQ438BOmBElG5wjuL2Aw8NMKWjG5wF+UZxSUxOagSZ8
WyKSTAoGEcywnQaUw5EKQ3MQJF8nSBxvi1xh7lDG/nUy984Fw3jraSLOE16d40IDADir/VvkVpmj
iZ+oLCDx5AzjQ6Z5zuhsRooxvjEnXmNQNFbat70ih+cx9kSkjf1UYBrIhJBVEmtDd8jygCzQw+3P
Er2pRVQVC3ARyrbwLaT4dCMqHYrCd4WIyEkRISWixILaHg/wH5Nh3JyYELuNCxEz2/3d1JdIZ/GD
F568eM+8vkc7ezRocp/jRFPlXg82VLjC91bwgeYlpNPV9GkfDXWofsWH8Vof4jieMDr4GbN3SgZV
T+1aosm69pG5JMOuh8YjmBS9U91lAM1oqQ8m//M/wnGsxQhKmiSHDSNGS+nKi+hbkWgqwUlPmqwI
ZvUgZkf2bDq4XyRf91GzVi92DHb7vSn2hJOvMUyGLE6c7eB40TDXGVUg6NGj7xutRPbzapaM/71g
Yue9ja3EvrGBAO+KIr6XBDPcosADyG8xkPDd1blGu7BkehI2ps6WS23aJXtFQg0LLBLZC6gU6tQr
a2IImzO+nUuYEUTzoz7CB97dC03cu0SmQuFJjWhO6+6ZCFmIT8jeltnpt3/U2IX7N7shT2M91JCA
qQVNAuE/7GifSXEkpalsi41HBDXCtyOyTVcwgO328yhFNc6VtTTF7F1W/bYiThcg0EbS/X9LloES
/BA//7Uu+5ETUEecA74rdXRh4/gnYS5zcPO3IaTZqsl+UTpGZZAiRf8DFQFLEuq008SqjfsVT8pD
33UL1awVxaOdOaJVil2V1d4QTUo/q/cvu5TZ793yE5Io6RpdTCl0Z08cbIwtu6dvPuvKrTbvaIP/
2LIhepEhaHwjE/WTUCv7QuV58Ta7TVSYGdidY9sCsSB2zLZWzdG5KjRbJRoD1GQsH1IE9l84bX8H
eCY9VNvH2LjK8OFPDxfGVEemCKOHtqBglswQic42JrnQEcsBQB14WJay0wjl1sh8zLbZuCM7vlYw
E9zznOVWrf0z8d1fS9ZdBP0SvGy/GHMtgT1BNCGn9K/eNG3VYgxDzu23MgW2BCiD9r3Bg2BjrPfP
j5scQQzRhiOP5pz1PZBdGJXAjA97Bbuut11ig6WsT/wLiSDqo9Oy+Et9R9k5pjiTl4ahBc2Bpf2g
FtQLxTWTbCxKhgtwZgFk8Z1kh9lS2TIMNtzW2e39gbqB7eX1hpXz+JqjQl/C5SssAbIKwLLhhMVL
7zL8hp7CrZrrDLr4tOQeQFXjYiKhJEcq7efAANg+UCNwZXSl4U31K6yB5sEaZ98yE+V4WRZ4Qt8X
88vqb2mm+N16GEKf2mV9A7IJDQWWVUP5uhTQA4+7Q1rc2sialO0u4C3CSyHSh6RkXCWuOTge/loF
5/xq3xBlUzeK4mDHnaDWEDNKaimJs0KW4Y9wkS2rN8+NW4Dx10BTCTUN2u5QVS+Vbzyby77SMHHI
qpnjWw5S8Ai5O41UcFsRUx0W7CSnU0WEJ5STVL/3hIgrInVl8XkbAsVgDCmGk/Ss8KrhK1nnt8Cn
ISMbSbOIctF67iQLK6iIN5K2TkBQkcBB/yU1eDLnUDCUXSFJIlZhJgsGUFl4/b5w0fYYb2EXbJ+r
DpnWE4PAq6nody57byiUke5zzDRwh1+x76s8ym/4bvWQWaZb/pyanC+Q0dYjk6ZSjgBXqDWKQfu1
ncMa1DF5xrxifoCfqLGmRFDnQsWWd659AAmFsRYjNLnTzqsPxRYCskqmMLmbg8LT7E9L6olzgKUW
s4tjGwpUGBPnwG9SvmQhgbIAbsnKvDVUO+g84HNwos8q7wD1s+b1hkR+wHQKaTo5RQyZtZYLN3r9
GSggWitcw4iWa+5MR/gdcM47a/yDS2BMHEtfPe+vVuLHtF07t7dsQCqAf8hRHyiRIVMmjvPv72jP
JXLVY9NcliCFs1FwdPss8E+rVAND3B4ggEYxbaJryDyta9birlZgSJP5T8Vz8mc46Al8yLG+4Mw2
3A1bzjLJo0YmXO/KgoX58ndQlWumNUWfmqSFWD+7uQktCEicD0PZz1jerquIOYfKRx/Xy4TUt9zm
Mg+3YL74GH0PFEJY2QdUMtKdfiBmF97cr7/KJvtC9N5+lrWR24PB1GI3lxL32eoPCQ6vx7qnlDfI
jWpFtprIGsLQ9CTALS57cgBtwECwooxeZdAAztrJw36h3K8eOws/TlZlPzNocbXzRt/Y9NydL9aJ
k+vBJ4XrcEr+CDoBBj0F1N34yGyQr86aSLuqk1nqwJGrVyIeTmvhga57ZfjEJ5rYgTfoJKTqAwIK
IU18djLxBcQdN2yA5FdVIckPjQLAMSsPq9wCWhQRDHs61rCBcdfBnvuwXxeBP91XccG9rxM6Z/Px
JtvGD4qy75M+m2eRMTnpNvTfOOo/UHX1C+ptZ7xBosmqwJ0DFKEZofAm7lA6WZOch1RyI3ZWGVge
OKaNhihQH5gWAT6B7B71IcwNhFbgaYh7o5wq/qXBBQ7BNeDwWgedWsjZloXrdFslr9APr94KntQJ
PjR33GMuYP4kSyezssUGXM2R0AXoIzHY6OfGtZosdQ91sPLWjyrHGuu/S6heNfGtUWwkZ6LVN7Vv
19RDJ1SWN61M2uPCGGpDRyKbgpNOxSBgGvJV3Gz4AEZhr5iue9UNdUGM17+ntJEFB7ZrNQVtq7T7
SBpaF+eG5SCDePFOXA7RzLeTFtLRtVac+vi21RQv1fxGV2zjLlo+HlQ632deI0yrfPazTOMOHQv6
xNgiqSV3iHQVLoet190lTHzkZ6yycTph7VsR7PnDd/Ove5QnV+C39KeZkpc8pcr9UwpmcxPzxd++
IARDkTOMwM5gK9gRbc6tsDF8DzOufMCko7cTvu/Z02pEWlZkYq1Inrsm04/WqD0Hhlq9ghmwpgSK
p6QgbHrDHQbzNWnx4sJCX7GB9Iz1EYXEm1oZlPUhn4fD+MzCTiQRFH61oVcDhrXYQcW/mAplBFyA
oduMQJFOcn4ll0xiHgOUMsmWE8YO/VkN1nS/zKid+wzknlFzES8SnoliuwBQ0jSWIMUEJRYFXmQ8
Ka4dRk+UB+qrCT5fYz7ersS6nL4/fxnEHMRRbmMFVrVvYzox5F/+8W0LrMUgNqAY9GElAh+Ky0BG
+2SKuJ3AviO2v2ppuebMswJr47slVUgzg70hcWJtTGHStNZmAv8jVibcuxYjko/3MLg8bK3d4Ip7
xgEUEdn/K/sztlriCHZE7KzxGoLYZa/knz5OgLNU+Q1Dl7a6V1+KtQZLHBvCsn8B7InWvBb9Nugb
HwAG7tercg5c2PcnVQ0Cv79TJpSrJVEQ47HgymxwcIQwpcitFtc15qsQJIZQlhyLr5Ay8+K+cPCV
YRroj/ok+JPLqQ0k8psVVfjHiwHRlSwk4KWjNXDEP7s9Pta07IcPkppp1toNf/dcpD1HgYP3ggbX
vatPolNEr7Jg6bETW9sXbMma/1aRFjgpTIK6j15C+4RLi37ofjFdwE2Q04QtZHqo9UfmDqgtC0Bm
+kFGZbDjy4YJLW7d/mplB146psThYDw8hsHrJo6xt1sfTXK0l0PxWxQmWCcEHf0mPG3+mWXQz609
G0BVeiW1LVywEyXdemIzUcKAh9K2obXOrrvWQp+gKUc2RAqGKlDQSAUuYnp1pXYP3xqqYZc1NZOK
i2Kxm7bL/ltKzX+KTmjT9KGcu4IRd5zIJRE4a2OdP2oOIZGHgFF71ValhU48b3sq25Qw01DExOOH
ngEolLqktoR8AeobxEfqIBIuCh92HL7+rybe413fvzRn7V7fSZxNG9t+4wToZwyzKwfQOxgMPm8L
K0NoC+Jc8cWeyogp+Q1h77oJbtZ40ZHAqcWHzmj+YjMXfUvWs/5gzeHJua7lVdoi9YkUd9471/NA
1qRqwN2NE4JH2bwN4N5RitA2tSxVfmDJj1C5hbV+LJ+Q6q/+4Bu7m2UbpN8QyeiURnYAjdOHSugd
inEa1myY0/d7IJ4FuK7D9YxYfXimXsAxGpoMQdjD1wNySGjSL9GuszGqAycmyjAtvzJIb3lHrwaX
6kZxKcj8rxbY4GjZoM0eS9ACj9w3QlX88MQdyWviIvd0C5slC/irmWJInEUyX1Ssb+KQgGBpKaAw
7H3nniiid8KXu940CmQl6w2+GgHA2hSQ+d+Bneqea8M5ytK3RIvOi7BZlbguy0wVOcjdSWOfLhq4
VynVwFxF/CyrduVEXQaeQMdnr2q6iHlzZoj2LV/vhc3EJI/BJIlDFPVaP/RwpqYuIaLJocvSPfS4
srdI0tYzsiXpyhEpi5qjLuw7z4HKRKpAQjt94JxX3o8lbgC+IUpWEsDR3IxvaKRPVvnLTBkIgkTj
uzk2xGE8ZuvNUmls3wdg1Z2+t1EX0T3x9tZDodr+K1fVJMKdi1ERKsjM/VJ/gk4XrZNCFz/e+f07
Ag6jus9ds7BzXdkD3sEjgZGmFRSFsNCxzLjglNUc6PqAPHOna3Xw814QvSstXZV47JGJHl9l1N76
DjigSrznF1YGVJiSE5tX8Ifi3EaAFU7nNN4WvMnYQRS6Rz++De+nMFDnAebotF/l+3IixaHEN90P
uXZju/Oamn2boBYYED4rch4AxjvT99PUJhi6ebvEUbPNqMEcpGoN0NXTh50k2es0+S805zXZ7mRe
QdFtbbWSuEZjGmS0GP28onMPYFwkFK9p2cF0ZKYdfx3yZZC6zWmb1WI6VGkNpNzMP+Jkcandt89x
wONcUDUobvws0WJvjyVNqxEXuNc3t22NLzUFLrdGXBBdsaO9O6njepSpsLfH2lkGonHSor/KVGba
wolTgVfFHT3/5L3END5Y0gUqrXJTsJ+JburEqqXwUdhzM8PnRIhoXzBxPax6Mz0iOUychMG+IxNl
2CNJba/VFLit1gSZy1khzu3tmKSHBpXpEwSvEK6UMYB0xq7W/1Co6dJF31tNOq5HV8i5s6XYljwh
NWkrMv9X9FgkxBaND6YHbVVdsUHRxm2ALUNx/gMAJOSDZGf8Ah4WeLlJNXcNzZLdOLELhFY3jPA+
bdZqX8i8AviKftWIW7aTXbK1tJC89ob8BpsiRC8exULm67R5NRXl+Arfe1GmmRG02DTwu3ycymQ5
OUsvNKZHmTwrXkcXQlFSBOhu4BDWd9KXecjmfA/sekquPPPs4KHPCW/kR30hqbQpNBXV4p9k35si
UU/evRjoVQ7UxFj5u9vAx9YfFE7z+s9ChR5RhazW3alYcPc/r21RkIda9RzQzFNA9jRhrh3Y24Qs
9itaFSjI2xb+HVkAQbMQ4W8BgE1WT575hhMqtoJj2N5Pt63syu94f4kVnk0pHnCy52Lt0as970SA
SXKKhSx95/ki1jWy723O5eU9Av2L0GsWb1MvMl59gun9hwvXZGS0jcBGyb9bBhEBW+hXdC6ouq6S
Juyf66ygv9MZ2PHNPtUHUYIQIqYUQOdOesbUgxQJfBf/K0TOCGNm6jf6A/H+jREpxrUUYVxSbJuc
2apF5Q2Hw0v/ML19ME0cTbKBwm+0wYbyakpXMp2D0d82lG+WyflK+nu9ZpXhnPPlCbxOoZKm+flN
8R4nEIZYX5UI+rIds885aodFZIHbMHzJc8tO6H7Sf5+3/lmgor5/cpLZPcua4HEzHn3sSbUlLuOE
OK6Nx3Y4nXljd08/0BO0usPUPZ3dn2XDiRcfZTonsKGAX++4UAY/x+MzX5atXlqiKbVII/hMImy3
s2UmfNBdU5RvAUwCJfouJBm/LiQSDb60T2yY/uHpVds9CxcNzu52BZig27ex/fSmwItQg/Pze73u
OxRZU2dMFsnRnZCYXZWbagh9EW9bEJmBkVnteS61cvilRjcSjj6lQaHiF50kACJYax2bzjJMPPXd
zqnQ8Fh5e21KfO5d7y0W/INInH4mPmwl04B56RAFNWfdcBoLV++XAg0OyhfWkiHP5bSor39VnJcu
Xf9V2QfR4/PX16LX1buddZZFI+ga+E+a90OyVGWEoPzedPWoYG2iOYqsVzKiOvLCP9UuIlQ4hhf8
EOHrsKC6TdqMoyiCpuGcSVp8wqACFqAw9/yrSiTYPZwiUNGobivjwo1hYYDf4Fdh/tSF4kX9mRkX
+NsLYYMG0iCfSp3z5C5KB3tB+83Y6ZUV/wuos6Z32it0bxf1/zRyuJNt6YwmqmHRXnNudAD4eK3s
lE36oiQ9ZLegoqSBdLg0GIwgvGFSwsk0duzUlf7p9Fi5rgq0etaZg/X37hAZmBuLpVmddILUnTBL
Cg/qjw9HP1OoVxFBLvuh+1iyyDIvQZa1G++0ygFGk+AaukmAEhL1KUEF5GoaoUPRni/q7UlwiB6d
1U+MXXif/TjujWXtUAb4q0NDNmj6ZYVD30uyyzj6lEhJKet4I1zmVLy0i8opnDl/mH5ODqdMMPoI
/AnvBqGh/bGhnBuyTEn7Qz0k0wZaVxoIevwmZLAXtIdXa0SyAns7LReJnHyfhLaoHOTwQx0baefY
3Y3pjblRip+u/5xWEjmEa4hG5LkHn80rHYCTJsTLIUVTbTirhyCTAxpFWteQLCI7YFHidim9RqP4
GlrT8kJ8k8k4v9qppbLGqfTkpSJwv/P3DwhYjdR3M7dWztfuINIORx8vFQlOirRyCeJ3XF+2g3E6
dn5+H7OoZiE+xhE9amQ6vnwCHATnRzZMfxectMmUI/ka3yMS6hRyqhWUzls926npVXge/i6ErjYC
ECCnMAeWsnLtwdXvaHLVPHXv00GTYlcTp0v7QsCpHcNg76amziB4FQtsmEzkCby/XtUfEejO0mJ6
pTCD2v/cN1qHc3ZzJiiW3W/dryiZwPeJ+onAC6fgJX41JbcgjR5hWv6fCuMWFw0v3SOR1wPWI1qO
tK7q2J0/R3TyUlJsImzo5nt/UvmCLa61YX1tEGpJmx8/jfHLKO7OiyJgfryfTNgYjARDSjrPcK9u
pUifzDfJMfp8BbQmNCBflpuav9SIEJ+mT8tYm6E1v+GP4vDyNHXFVns7jBbLQd8ZKWhcYOyI0ImD
V5Koomb8+B5S174de90GGlXYwl1aV6zuXTpWnvC5eDfReSuQZHx4o9bmvA7C8cFvn2YfoudIhhhT
S8BtdAWgXnswJYEbCxej6rK0SJUNR6qDLWqBq74nGkVNYYM0cDviSdXMmEDx1hmBOTomK/33Of5W
Jb5LipHbI/dRpFgPIEfHnZjI7hRDCKq9eta20mcBFjVxFaesZXtmgsX3VTvz+aIhtKzpwCNAaZ4t
UUxKJUrXzynIJTZROk3GzKR6cYaF8CogFdScc95BKmE+tYOw1J5+ITU1coKjZ6NqJ3HrUzUmC0gv
ylYR5oXh7blncr37JFKAJnn1cdEwQUez0fcmMP7j7ySna7TdgtyHYkOSD1mcH8OJrMGHO00u+J/5
Mtjd5SvPZP+FW0ZBkcqg3KpSRzcarFqXqIroCJGQpmPLryKXz3ObBbJitACILBrXqXINc/r7suZe
bAFj/F9VHNuzOR8uHBcYyfRyqHNY0BcDFVso/4d82g9zoG1fBI23th4wYIHep26hCECxoWSL+WBk
w+d3NZBWGgFMLwnf0nDmHOeOGk5HoXViIp4dWjltcHafQ8Yf2IRNr31q+TBGJ38KlWMD0FSqyMhX
RMXU3yFL8eY/bwJkfcQojAbxWjWFiUj9l8PD8iMBX/8Zop4/l5QgTikC4bkPDiZxvWTcXgPx0rCJ
s6HqGoiXstU3K9qDNIGRU3o4wnBTN03hGuthi0a5x4+aDXcJA5hszGqaxzAzFzaH7hohkNPMdNbM
Hgs8+w0OSXb8W1K2RFVBt29zcNPoxJHuP/lvgNvUH3Xmg8sI+qRrIoVhC7fRYZ7ITC8VHiQGvfJ8
ymUUnh3txeg7OXYTrlLVO+IJ0NFMWIVm3LPxtyfJf4ceW+VLypXw42VKHUB3wr53kKIhJEPy7l5o
uQUVRgKGP94BFgZaygy3QdHfuzun/+NXP00+lzlOMIspg1aMm+0OY7qUvffBgFNfYzXqsclWUHJu
FpQ3VV0S6ng4d+R86dqKKGMAJ4Xf69ziTjtL9VL8zsDVkqPvC+KDB0MMt5/C0530qbaYaUR85a5W
DFl1sciaDoYlpcmnFnabsU6Ou4UmbfyFzRipRxxfXeLfgUVfpuEWOuBP4H1G3zFxki3nCnPnSBk2
5khYEdZ4cBNBZOPPHfXjXMGkyLAmlUT00CTaeSA7FR1qrwUoYrsjPKSNlKoZvrFvnSaFrwJ73S4+
kYCuPyByy4SYoO3kHa1NyUoIBV7jbuFI15xanjwEPMXx4dd2vZBur9S9+/LbS59pio2UzADWhCRn
snwwFRTpuHgkazJQSS03dQcTs8qK9pz7iVM3lQ/1npJ9sVPjF7qTqjwspoH17fsutWk6TXlyLCC8
VFL5HnIluxH7/NNpC2oQM2qlLztO3ZFcEfuy7h5JblXBLuifHpxgZIEfj9+eyt4p0SVNdwHQ9J+M
Ivz2FwYccSdgz06UFHMIPAgjEd+bKfekMUXY88MFpe/UC/+mBdT7Y+Uy8ZPG1IHmRc9wJ7IQ9Pma
6yab3gV6Q+xLHzxQ5G1T+9Umki6qLnZogJMAZQqRR+F0H5OCp3GSQvmRPmsyH/4Nm9IdlLO3mmWk
oNYcMQADEdNOXmhmqvMbK80FLhoE2g5wZJq6t6/4aMCbflyONvT7oFOJH1nl1rrhatbAIlgeJUxO
vtvfkskIn1eZ2cI5+ZhKLvKvXIx/fQ0DEqpIjLjnoAxpBn+O0h4Fq5VUU9+OJF9Chbo/+wkBMXlp
Xj1mIiPPmBIhWk4h1TFlFCbeFRTjptrsa5n6gQr7j+buZ6O7s3nvdG2gxapo2JIlOjN5QmMY4igG
3nIlwdjeZuTlcYx1VjjG+oU4wpCjKNzE669WsRhzJEk7x6EPVS61nZJ3DerCONkdMvOAaXP/+ICt
p6wwt6xFqK8qZnDQ5QQLassyaNOvurTM7gQ048xce3LmYbFo/VM5kCmy50u9z3X8ZKajnMpi8N9f
wt8iYKCgvstWUgG4xs9o+Psesunu+yP21UPM59J991ZmzAKcOKua4H3H0u0jiD93oHMl7yXJ29fR
0/ffPJ4bswOduX66iJyZUykN+ouj5gvMX9AUAXx/htUFOdileXSBiVGN9Jt+tXp27HdUJu8UBGj5
ymE/OPTAmu/jAf+oZsTfZ5qQa33x/YmzwwipIW4cpcWP497+cMNy4K6ON/O6zYPnXwwM39UAdEbX
0FZjWBMfLMO5/ny/DtoSib6ilCpkcptX3itlMypW45LU1WKUCVr+ShVl6pSiUDWnL5JiSAV4DBOB
weZkbvp2aQZQUtJvyYQ5UCUjuTN6cfvScTwt4+sWYxKo+SD54O78DdN/2zg+QUpGYtC28oXEq3Vp
Fcg2wUomxasvqZ1+8WuXdha9Zl+PPcfkS0TAJyV8V3nOdd8xGqLqgj6iX824JINQNyfnOEopSwQC
5VxAcPyTAe4aUxvI4x9+O5vbcFsMk9dZmmy2T29LajVIhpfyA/yPNTCnm/Cq1r/dSdqW3jBQVL15
G8HvCpm7WnVNIPtOCmIdfNFJalk8D9NFgpZYhd+COm5UZkFDlv9qMTYZFc5LlhsdxgtvgpYYL9eZ
IAfcV6ICY7ky7l0XRvacj95SaRQzNkEsndotgTj2xtTxE+sAoawifOWhXj8B7BF80ARycbLXsbgZ
6F9mpuhsQFXtId2X2DLtYpWwqwlgY4Gh9yt+gmRXFZmiv6fB6hj7oKkPitA10e1pEHOD4PaChdtp
ajRBdDi8q0t8QFoDifx76CMtjQsSvqXto/Go89e5qJtMob/9VYG/SNrfXnopovjzM6CYr5YHt9mY
RTfqzozbM3JIKZnM6kpM/S2KoImVAAwq7+0AY43Y0ofk1NPhbi+0HSXMNIv7vvG1hXu/0G85Xc9w
RuPda6vsbbfXQgB4pPbnk6juuJsNWi9+/cSOmIdZaVoOXRWC7hNE1HxtTU5fzUH0G4RvUS2sVELI
maPF8XH9gM6Sp/JSk7UfHpVaxVogztCH26U6fjcG7pTzlDIn+l8bIuoG9dxWXN+QD+Kfwrm00jMl
5KBEWtPXDCCX0J/GW4iLG5KIJ8pY0/VNCoSUzfn5JTjv95V0Aoa1aFXe28DsZ0qrmCekUkMGdoKs
9KrIDr/lAgi7K0JZfyXx8mhnwOvgoHZFaG+X8OWSRYVtvGeGTTO7dsG8nHYcaR0mtsTa9bzraKdZ
RX3wQd4wuw15pcaYG3wbEardDtASyEcW845wwNsc2fb/bhxY76Y/TdSU5OUe1tKpr1TCIlY6UQR2
m4lb1sreXx0OVFgCcZsDRbjrFxqp5esky9lrQIJAjL9h/CrCWsVbJAvfF3NnS73GwKGZPd3uPTOI
KQRqK5Af1E9qRV8hSX7DUQ7JlzRvEy6t+sYeszPl9DuSHGx9z//Z0bDFYRKZBqtPBiQjdeTUYSdx
9c0ifYHWRZ3HrbIBtjVSmmBytKgU/HyFUIx8f0O8bN2QJNXBlGf3UKly/puY+4rdKW3p0/QVdaj0
PmgJP3lxgksxiFc+kBzCPOPES4oQcM1K+zP7L+Kv+zrsxi3legQPG77vftBd2wZh/Wvxs2FOp/Ra
dXGp8/zaGlSUzQ6qF5gaoASfpG41GJfcdOvx+grL1a3pOnBoRwJlkN9vL2+d8Ol/jYNI1RNv72P5
byx9gxuutyfrSxosWi6Ij3te0vUd4T2T9EX3kepXJdR4hRVDof6BR+7GAQD+OzikhswZDOf62aq8
NP8k8MGXAFOvHTldT90bFSOkWDiSTiC1+01+CFCK0Cm/RxM4hgMQ5USEERimOeOqLvrgZ8FqnoFv
iK/JUE+xny7wvBVdkAASHTCDNThQl7pFxakdpjoMCLlOFqlEl/x9nZ7DX10piz028B7dSH3vAmSN
ltX1Eyt04pizpdelbgvKFodmk9xCQ8SzzJ+5oyMpkrxfTWuVrkRL8tkiz7XrFQqzNkJ5lNAdFb6P
x/I8VOMTxMnJC0u1BDavAoglEdxNlYGqbDVudtlnR3MAbMTFPLt4+1Emzkes07eJ2+wCGulrQlbk
lZXZV/9Jsk/SLfitvbE9ItvKUTeTVPxge49nv5AvJlMErIV2/ud+ANMhuhgLYiGaIjIRq2PMIN0R
K0FFEt/a0m4EKn+KDrLMnrbovvrnL9pf04wR3C3rAU7pC90YmEqav5HptMn+swq4gpN2r8oIrNln
l3MUr7Bo+6+krwl/FkMUJ4PCgTezblrcf0QrVFJBjULBpzCBRh818w+PAOAIqTF/btKiN71JIWYG
TjdMkoj7dBd18oZaqXAsJKq0B3KdKT6PbzMYoMVVgtukeEzzTercVdH/Wdez4SDrlXBO0Ig+tov+
8JVVatjv6zkzeDlyxH4j1Ir0KiUHJZGRWoRNfVE6+mKe8DZXdhTZCBgaZr7hB8nu50AUt313zxPe
C+Lk8EuTDt6mdU/WbAKUEC6hCsj/1JuzmkHgBN2CHpxvzqq/D/0lXoWrN/KMQS+n0yOf6MfLaiBl
ix5UJZoKhdQiw1N6q21N3M3zWh9kTVN63UHYCTQ7EzlrH3BuBypIBt4s8Mc6VyYq0QuKLMAFnh70
hbHXE8Jyjs85EXIyAsq6YCPoKWdrJ4PFp+Xed1G+007J4t7L9gtrDAhh+6gXRG8NpO0QFi9Tb0gu
XAHCd9e34belf9n8E8b6KDGd8QfEvAL31k+/wT2MppJoOGNZll/OsjsiiNKvRIDnFwW0+5tyDUL1
JmKLRwDzsrJVfZn6A1jS1CuEHtw9Bif86SCrE8THoNUKBohKcVtXLUE6pcb08koD7IYQLph2h7cy
DuTsFEu+ITs0+b0U63EcfXquTdxEUlGVn6HXs4esvcWVaYVrpebUOJ6Vw0wuV4g6uVLBca+t3XJt
37JlePPy4QenMQK+lxdYgOy0caf6tMBh8Wf3izY9XncMq5tzkHaGbmHled5SCDpCbwsJwcM6wUpM
SyKFdaz1hTa/qp4Q7SLbgSm1oKIgjR7U6TZTQNVMUUlEBDBB+TCSYN/sSgV4Ty7WhpUT4Icdevoe
xN8AWCOHKvIAE102Ws/IYB7Zuzm7v4pixziGGpIPiUr5/OFH8uC2EdoAtWzqd8RMP4j3AdH1EdqZ
lxY746GN25ygqouS92eNqTxy4nluJLXY2B6plp4nJo+Nuzi2GMmiB8KQS4N04iF+i+zsS/qU4KZB
8KC4sHQ+SGcVvDlhb5Oq8nyPcpXNYtKjqVk3X3PhFlqtCdPUsuvdvG9ggpDwtKUR5SuKzagrOwbv
IC5xTPR+742BA/0VD5o6NqFVba4AOq6G4eOTF2YGD2MzEPwW2Jtgl5E4GUd0dSUbgy1a9z9tMV7I
08ESS1gVQ4ISL/oXdt3RkhIH2pquM2to0MNkYsyhLNh2w9RwIyBteQ6BPgcPazNUkd1fjHhHY/m1
pU2st06ApkCu8lyKmPTGutQXgMm2z/UKmtdrf+2qTW+PhEBNKNEW10APYOVamyBGXWi0MV7u4IhC
u/wxzwb/mKh23J6Hv9ROBHBf/VNWZUuWhT+jnpPYtemhLhpmp5A9MBJlCqfEHSlCdfhFsCkAFcL0
qgWgi/X9Han0uSuZgeq9WQYdMCJ1OOzXB62cljXjnw+N2cZW2W92i1tqvwi7EGYgReu/Fa2V7XHi
Lrz/IP5yDcPDEMTmzpWFwjAnBV+uPyeJwsI9WeFchC2ClyaXJDbPhf+qazHDp0Nsrr33lolvlIYG
euF4JjrfDP50hvjhOnzoVij8nBw08gn02J5RvUeaUXc9dtJmEphS0BoHCxnTOUitxNPN/WP9nPMQ
1MPNhLGMDgjGyp+/uMiMS1o4tudXS4z4+YQaV6HTz9DXeq4KfbCFm7JZAdx/W0Ezq5ZcfBgovUTn
M5JspqvH6K0n9ES/GccdlrUjkkpR2FgR148IuQBiJqZnDPQCof6glZV0+VglBG+zR9Fr3AvCgtM3
A2ufZCStwwG5IkQn1AuUtv9B/6lk1VytjLR4xiBv18dvULdy7vzG33Jdp1RlcdjuZRy5tOZAFKX3
60CavJzhMKYz8lgK6nH6tKJfTM6yKUX38FizXGWtRF9RCcrQNFk2M6auGwU9kJZCkzHL71OEQlIx
0q/Gr0AELyuhPgEtD4kaC5Ug4HS5MWqpN4TzbWqCbkKjPOd5XXwy5IlFp9t6gLVQd/gSN6zw5XnH
0VcpVzXh6BzoUL7ICVA/3ZJvA+pFGfuywGDsLVGnSSLTpaTAuaKzRp5rB858FmJbXrUakJNwFBqX
EvDcN6zMAPj5sI5wlxTctlHa1Ru8Q+ThZs+60OUhFlu8GTNQv0YBNFs0Zt6RPEsMVmANstv+j3Yl
Z/gqTzBz1IAfT95nloCap9kQ+7jfNkI6ZKFmAlOQzuT0IRObecFk77j6hE5okLQZCEt4WH7HXmnb
ncFsBMhSvk9hWxfozHl6xeD0JlfQXbw+ZYLFHpLcm6jazCVkbwmNYcIDo1JsAzpPbk8ypyj06e6K
ZgeMHsyCCVrVHWAQ/3wx3RrHxyZFo3A0jUmdDRNlUXSdqzA/Os/pZGL16ohI3Kvw5qsuW4933H7s
NURc2B37lMRLhZWxkVB0xoUbpKlKiNWi6Mj8R4VIIDM/qvWJH4XzqoRTHM2nDeyS3G4aoyXR/MGM
gjRMGszsstJpQDvnZdtB130h+crm6bvboPVSFywJC2eTz9JyYg7W1BYNK5F96gEOXduI4eqauFp6
Pua3H9R85wz4e62syCxRQeALULGlDj1qmayyWJXzOSN1u98qW5oR0G3LhXyx/oFfW47zTuxsVF17
YJZWTXXrY8GNff/J2QQugnUKBCbFQG7WgvBcxmEgodJkvvsy3hB/dQ6/iSToZhYWMyqpQ3q7gQIA
SbSmM//ZcEytMNU7jkbmsatGneaurMrDGa4EuKwh+b9dMAoOQz1Ppc2uo9TM2cl8IjMIHy4rRvqf
cY2+sbpTB+LLwLSy78OMXgJ6roKfftrrvscOwGK+4oBDBr0H4D8ulhul58Q57L9tURzNmlxZzDnL
QT/31kjLxyPAyCrEl7W8e8a176BAKFUcCCsYpI6PN0ITDIq/MZf9b8SwYl9rn2R3sjo5N1J+cPT4
qls/pgoVbgU47dTkiQ1TtORT+zFl61arEFBkebpCDeef6hzSgctwusa2M4KuNCgADcc8asr6wTwK
TCvoRPVYxpRpAlzwoWOE4EY74u1USN1kQ87MPOuj8Dnt48iuKVEJ5qzVmIWoqC1tTVOu3QzESBG6
Yar6qz1LvonYAgtrcIUJRENpA4gj4r+aPU+M1bMrh1tD+yl9/B11cdmmV7vwRBWAOBbzFsgP7U0A
EL42oGf7e7Nq/c4S951FAjSS68dolkYFf392hSM36Hep7djP45f1VFjtAAbRCBsAkSpBIqy0tOMz
RSm3ChVBPvD7yvps7S4DCWUcsrfcm++23MMVcz72hMdBqyFs1+9YHR3ZgJDdND0Jo0oC70z1H9Bx
UoupRXO+KnKug2S38u3BwwakexpsJuJJ4jizV+ReV6xHIaHImfTvDbcClvZ0OC3yWvK9zzfyp0HL
MQGwUT321Y3nFJmlf/JInlfRFBA4aSuMmbzRLKmPOSdFY2EwuHyRfarFYa2/BWHaZR3ShSsS56p+
Dp+MdOtfIR9PHN0klVH9gQwm4r/LpqC77piFw1rsny7hSRwqBsEJCFV3KWoROJyiayFYqnXJVLtD
tR9dq3OItVPDxKgpYF02+f75yhwVbW9hGMP9ajFyPxH+Q5pPYQLYD0YLe/khEXXnxGjSUY9xIdNJ
oLUe6FlJ1GfYSvvNQnKtGVqzF/EbUcs98+MsW22rMbMeavIqRCoG3C9vSVjtAuoHGDa17D0/ojS7
yvv1EsN78rQTY27t30bU+T86aoGlX4s7ffBMdpZGyVFHSMB7m6PvaBLHemoG+j/tjxM0qc46B6V+
Jm9KYZVYugm4lpxPFQigJdEbp8p/FIuN1rtxYi5RI+UO0Wq/wyNC/gntFBoiLDOxaI+eHRBHkAqI
OfMblgulj5+JlhBpIsF65H8ONZg/viRk9Coox3pB9kQr4aPQCJpeswdTmejtmNsWfZ/UGSaDhVQx
XnrK7xZojR8fFeltHrIEqsuS8pSIlgqajuDOswaz4aq2mhJF/0IAftcDx3HvedLnlRhyc/y4Y5hx
K8EI2tZKUVd0BkpF3IU5wBJZpDv2jxF+J2nXzrUSBW+CXVyM520djqyg60rD3fdOKpcUHOrG52E2
1Sr4hhoH38aw9AGmkdTOv/vILav8sZOLdZKM73F87BxxS+UXZWNMXXji5bGUsxYAhcTXwp3P12UT
aOF/8n5GuChK7+EBD6dfhc+qXWFBCGYk6aM8eaSeY+Ijg+F/9rM/MSbmdDC6KuIAUa39riPCMl2m
pyzneSFFhURXLSwY45ysSaoOFcSfuNdCj6awunVP3/eV8b0TN3f/r2FH0RfGm690DoAXmpQyXCvD
PoT5VPXxSNzv5V0AwiEQwPopj5KpGuOpVKb/iOCV5bN6G4I7sRh/7xzFkHdBXUYtiaLPeAHip75G
mrQL5F0Fzt2rs0QddRrxPS5GTvsLKUOpN+Zt4x+HZWHH+/57nGIyV+h0rp8t5SiW1NQ8VwSOcM7i
Ke5QvGbFmM2XxfqrorrDnDvpQeHes9FKo6jTHWneyznQIXF4DlmvTCLRtRX97kNxeLxFbvOvD3q2
2jgQ6zbSScXGP10oYOy/imhaDQ3QbWvOiqEcGfqdpBB8jkPyvLs8vWH/JwXDqYM5XP/JIowV5RsO
c+Tx+Dz/FlSsA+dYCeTMZOGGn/JY78vw/MCE+avoXEtjgyVeCTiz+kV8G+pc5/p50y7trIiVL21f
1bhZMQV+9CVGe7/LDE1A3v+AHH2VJbxUoCyGAfbPZ/aZ0FHGaNK45ECiQQbIwRRO+xfvcwwkbk3k
jyntPZUJ2ZOKqzglLHQdEOX4nqREaW2TjAWuvFDLwQA5FjNUNA8jueYJ8Zdjv63EcyIfew3jreRs
931k62NB5yXK4T/rsj5UaSHM6uRINMnOeC/LsI7yIgUcgD6LQOyi3Jwn5mc0fYRaIjYvOmR6YfFS
APc4dxvhAh/iBOsedU7qCz0WNFXIqkw8XK2DRiuZELr13JX5LnSS2IDPgpF/vo7reUW4oImqAHbr
MqzpR2eEEfzP0LwMnHoYh+BNP93zu+7jUCuhVYF5z5w7TqTAom5rMGKccqDuiVuk4Ayl4DjOv9Fu
OyJupO8lRNm/l49tH8Qfl63s7Q9knsGJa6dmZY0qySIVrw4vdE6pyUWSHHlv0X3fOZ1K9bMPGOEL
aCVTcqWUx1cknC3IwobvHBNcDaMGqGGVY0Kg+PLIxrUI32yk7yWVmvM4HfKgnwSKPLSzg8atfWe+
8AzeSD6o5s9JzjHKk31CO3KClxzCOlx/QsseRvuPCI30lcTyfninhUwirf+3b7nQEk97gd/8hv5F
6sQDXEXU91vg6rLJEQHRVK7eeObD7tDc+LbnAt4jya10RjChPltravSemKxff/ftuU9Dj+uxqjPE
dU/12UzBNYn5bXvjJwdfEwsdf9Z68YvRqsjExHC5kMb9NPTu8yGIwl3EfTQRIqwYmhaiOkTO2OeJ
Tufj3kfa4QRjMaJU+DGfgiTKhHzA+FIwGfYsIDtcSQVxTwx7KzRyaJIJF8JcMcdcz5+86BjbRJAy
RpJ6bmyPHwI6RLkk/AL32cYSAAHI9tczofmKvPHLpDM2XywFlF4F2Cs8FjkSfsMKY4fBdmy+ID8G
SDoy2wClKDwnPegEl2jN/MZNnjt522FeWsgux9KXc8tptxRnvLkRjkUQvO14fQXDPRm4lDm0rAeB
kkDT1EdVyXVDsAf/kjJraY7oBmCGDQZftPwxbd0gI++Okm3DxjqqRy9z/Zve/+76H+4/Tq0QHvfh
gJHxGQHSzhCdqs/pz4mO0HTdD1PcWMFoP64agomVxiScvwg0kEZXBxG0HWvpQG4AzKm1DrSzzncA
b2xqfqBRRRDPwFpVR0gtRv48nDgGHsRHAquWYrJE6QwbZLwi2IvtSvBhqlNX4nHxeikgoZpH/+oL
g+O4f6ABgkwm43B5e4rs6Kv936S0B0eZILJ2rbeQ4pLJTEh1zZ2t9qZ9lph6xRYeE6gvsURFRV5w
P0g/AtMygoTEZ5YwFBdTNKSRiJlZE5gMDyAs4y4lBBcAEUF+V1pnFbe3oMLgeKY+FfplpTNxaq2D
nfxeBTMd7IzIgboBzP8c0HraIQIGB7F8rTc4lKS1WQ2IM43t4cWHLn55UcDE46nG2g/l9N7CnFtv
3CsVYhcS73X6x47V7Iu1TZS/dAZX/lnEKsWEhdKBzMSRFcLsaovQERLRtC3CpLHcQ43nJWopUqIv
PcXBVyVMEvsJbFCd+jMxNPsMwqDNm59Rikzq3tWHTMJ8q75KRor1nRe3qiTPrFgJATuJdID+KCML
70JmMo1gqdEFp29I7R0PUrkSRTXl5SKKj1glWZoGNf7qbNfxHZimdO0y6UnGmlSGtK6nXO/vF13E
KvZVMjlADBBWyZL6ORTRd+58793ndqrWGaeHUFR4J1yzkPCuDXxqtcs3CdFRuAWh0Ve+3mUiPVPs
/PcdX0b3yB5rSF86f++9u9typ709EubtumeeUcaf7tfLzgIdHSNiWWWSYQI1XuFfQV91ku7shOe4
36tA6YU7WN+yHEfzGBH9f61zhaVB5GI1ER40Y2hbQ+fL9kCHAbZUQQiG9ImLJ2a7qiqIsv+tp307
LqEfzRXRmq7fkxKk9clSFxybI2+iQKPF2X5J5sOyeg0LsIaHggpA2Ql8hg174N7rIvRQHbzNQYMR
EASFNLjJqyjqaM/7tiPF2fKhIirA9dnN/ICSXb+Ru7KaH4JVyOYBnQAcq0WE+/DmfS4fRcWlVIoP
p3YhYNjoAAzQeycUosreAcl1/WA5YBACE2dqIGs+7Iu84GXW4P6hApuY0Scsdq74OgWGvPMCNfOW
r1PMado0fSV3GgL7kmjlNjHZDP4TaVrky27dxJ4OGLJJf9lJ66bGqBAhZBJ9O2Fo5sDPyl7V7u5I
wa8xsLneSdVd8RkZXOp07+P99uZ3OuhWFupgLzXBu0iGkwXsBDEwzwFqLCc395a1OU75sUQ2jYMV
Uv6+Ab5qhm2lteEOiebYW2AVg95cleCbegWTGZNPaHwTh3RMTGEtYGfiW8Z+Dr+HJwlyFABUKlyK
YRxoaXsFM619saF37OALZbIwLCLBQiBYIAMTxGWEGR3X3TNbs9eyyUkoESbcgVj349WmOcURxugT
s/L9+rB66n5fdq+nwfFlWY384oOClapdQ29phjn4n7W7b2PkgJJfvlcJQtxnn1xOiNrt3a1TXsv+
QiBRyk0BE2MZ5RiHZdEZyov9pClKctxmcnVacLcXij8oe4zVa1c3DMAmIhqJpRt4KVfC6/XnpQYK
UIj6D5GZ7ab1G5ACUiCPboi8zhFGzFruR2mLKif3aiJ5xTBEjOauOSMuGYMgzuJJPRGcALITxhTY
oJ4aNbW+Xt4doPt1armRstfXReGLmpws61vvqB3Je7Ps6o5fHroxdvDndX9hivTzORkCdaPX2Y0K
FK0I3UXz275Aetvm2M+GCuziBmUJt57XeqLVfiP1W/3rGLXBOtu6b7K2Y/4fNtqU53fbWaVJgN+v
bWhVPOVrtqTN0W28ILHKd6iJ65Z5uesGPgqUqWUa3TU3+CsnHv35NrBXF0Oa7Zd79dEgqFyml3zP
K6zOvKoOhm8P01h9V7fDQnGsDw2Ht/EO6FfUx88p1Ce7OKO8UpJjHGj0cZIIx8l+3lftnLWl23F3
yjl8sDBMz9VMQ1XuKdY4kyYMce/AtZRSNhT5o+nRo4J362Yl6SrNMzPXCA5v+Iz0bh9gnr6Zw2vR
nXBAN3EtY3WS5i5TeLCxBLbsDcuYwi2Pz0iYqMqdv6v2nluZt6lPx/yleLTTg3zwRy5Be28vSawv
jVNj/8+xFI9Te48qUeQHMtVj0fTa4a6U7XjeJZxacPRb92tTLIyeJhRyTUmkDZx06NkrCTLYd3Yp
Snnln/dRmDsizZckN4E/j6b1f0ncrPjxGp9zPZaM3LlPKEf7LMpDimcyzLoj1c4q9a8iUXhNUuek
gWU3dQYq95ggbKtNu9MCi64JQoNbfC2NvAwqoLD4RzhXy798+GM0MWL9U+4qvU3V6nrL/zmK9wyq
oZX8ZV13NQ8I5rW6cDlFAQCKyfEZmHfAONDKQxnNH4DrEYQytrvBCMlXvZJh+FL0aTeI8c04Ev6n
gEm3oK4PLEphOk1Q8sJgWGXgDs1R1dIHaBcV2trE4Go2oz8sMG0buo3ji0xDzjvn0BVPDQCIDaez
T7UUaQvJR4aWm6q0wwqt1xQjtlDLOklGkkvXhLhmdy2wg7VMaPXGGvd9yTdPpevkWQrdL9E7lvbR
6PQa0zd7zRKtAAlEhHOOzpenX9LfG+WbWGRhyWMwl6qdKGyY/bE38Y6W1CG7ebbezYMPh59ALxZK
glmfAA20FpMKJkaBO0QSRx4kSigK6GsMTgDAWzvSU6QUAQuF9qMyehKGuUMMyIZJgBUPfZ4L6DQj
7VtuZWLWg22wVGspFk8Ooi5QAPWAFmDvSSIl2Yhjlv0JnBuvFpO0KeFj8bsTp96k4AtSyT+/wlC5
m1ro33Ku7w0RjGZwuSGTIoPQx7+H6+24ZeDde7HHEyvhs+0PVpBUq2e9FBRRzK2r2cDOGKmm47St
VtdFCRL/AmweCXjZMcISYmYKotDBIB++cppwzPEK+2eZGuAYaxc5yaU0GlhFsIo7imF5JBuhF8/l
KaVu0HZlagpK9DxPwdKcNl4aJotzu/9j1rEwvF2nY9rcbJp7smyw6cbqbaxw3v6kJlEXxdltMPgH
X0l32THuEm8r68iN+tcYvO+nxYbVIOLDV+SLANIoX4gGITn+1qjTQyXVYMG4E5xjbs6IItn/+LD4
nczEZIPqISCVRRJa1c1/4j87fKWMATmH0JE7s9RnD94GHonYXXV6YKFj1/T+RcurG5TOVljZCfp6
u+GFAx7uyjhCpywxnb1hWmpqBIcCr0x++IBIdT+RU/tL1unTQwvazgHv0gb7EQvbIA6dDud0sAj9
YBwO60Ly8A7NxoEZA/H4J+qKKhYPZ9ssXDDdvELOMi2jIOwz8qwHZSsFBsKhcF0ro66Yhb4voZq7
6YFBs7x12TGW0132Ya/ipfWjzi8TdL2fVHF1p1Gd4TwSWM2YismOiCcNCkHqK8V+bRgX0v1IXh3u
++YOsDin4TL9sAhlqUd1z3SWbVRXt8eJiDrdsENk8uZh3bUIWabzLGWjqwaonSYY6cv4B3BP9joJ
FPxfJfslzWWJaREoR06G1zj/z3dB72vO1emRu7pKG1tQvZ911HLuepdtMRZkIHaGOiQaP52ktYds
s2jPwn611FOidqb93G8EGdwNPOpdjP8SDpdEOD7NMrfv0nSlMKwsg2P/WP+8FOOBgrFinXjOJFyB
0y4SNo5inwW+16liHUgDrlvxyrLyjmvQNLqHn0mfRz7AdKU7CUQ9rJg9PoBFWOPmPU4qMq2e0t9B
CzR0gHrnqDzKpBBf0MaAvzuDRAj/++CyvcuZBG7JjkvfgAWqVo3kXwiUJB9ZahZIErHjsCrxagja
f6qkooMXTSwhAzZaQC9mj0d/Wot67/NO3BcvcTUIp6Vnq8Dz27klaEuvv4oILwfNjZAQae6icSsD
42PKXvVsHaxsVqtULmhJGkv0LHr6hZd0r384w90Grtz/k29mArLT5xyVPznpX3u359xV0LxCt/Cj
ODXNpWZ37qqlU+f/ui05DTs9VHNWoI8WgH0DA7V95qK0yJCmroOJJDuG2/dgSOf+/wuvIk3HovhP
Omdz2joT+x5Jow7j9o29IlT4gLMMCAHEOHdIffo9plKE7jcsmbDxzDKOr5wGnu6Y16dE5NqEXrFY
4wkkN+S1sUhAjlGtjgq1sycuf0t1/BMtyK6REG3z7jjx04n6PwzV6HmOiGqG2AVFo3kD2wvZ60M7
7inUG6QThpk+JOLivXvSKTG/Uok/kxLZeQy+/P01ZQ9Aqrco5FMgy9THWixhCiGkyTth2CEKzqmU
vFr2i9ObPeilLB64G2c4qqOMy7Hm2No8NsyLW8JYMCjSx/VwRMgh4tSFYyATJYrmDnn0vcEy49BQ
f71ZPqOoYZnFGS8yfdTFEi3C0T0LIfYoVwmWzQXUUJYMOIQ6wT70Y0UU8esPnsoHp0ru0sNFHKr5
IFBl4xmXL1+ckTS1yUW4+2WlYafd64YBqlQ31ysyKhELE33VW+uplvp4O8G1yHOHV5Oj3nQATkDF
ItRa2itj/eG30qBV6ygX45YIiRrsWFSpYGxk0BOip5Ap5svgZkteMyeDPJjhAfOTOpKzVEH+Ii7j
AmR0RgWGgTd9SWbJUSJHV+l6kf0GYfOUFri3QR1dAQcXzen6Bo9XihfcoRFQLcJwtfm66qKy8bEl
7DojPcd74bjGHUntntt/XYVSgb+FUAow22CL7Zes64rkVnl9NXMxewUzVXGfO6JoO+7MWyYsxU30
68C2PNlGa7XSuSpqQWUf6YRq2C9jkjJ+pYjraq4E0+rzVAzQXjVjtk+LG1msFTEvUBEzgpRjIPlY
+NXOHfgGquNru03uthtZGYp6mTx0wjx5epAmuNMeLLvAPoAX8WTXMgkj+XHIIJoCzlI9GYpZiD7N
7/D+GmDMbrqGpuSzRiKqUdlkZ/iz4RFr9DBFJ1YNcgcfK5a3ctGch0n9dV+WT6/gbOqyqwdbtK5i
WUKM9jcAGsXYZZC+zE7gjCjkkBl/xI5F+T9Wv2hzkIN6aaeHl87H22bYkj5mOUkkILXEsNGJ10BF
O/rf2of3EVBVvDFzd2g4Sgn1QDG0GKJvJ5N51dhAJdbzofQnBpm+laTTGQEgEQoM7cIHhwVzY1qm
hWakgv+yHJUoqI+PxfPASQYVR7/DIApzuTti4kT47Jk7keoV7oGEI3c8520iHnmbQII/d7ZJVTPj
kFkwLQ6D48YGAP1YKJ0sZaSh5Go/acf97TY+yRiRofGMd77xx/IeLa1j+YymGPcUkkngVy6peVFV
rjj+A/kqZfDksl+theE8B9yOSx8BBaBEWtvNAxQraU2aC+028BUFXTFwzSVBziqS4K9QtmXmdD9P
liqMqiZ+poP09qPKIBFVzTeUK3p0K8VAbspPZC/WvOiSw7muWNnjYczxJI8fLqe5XoolgJpDqUpe
D2P/wTfdKQ+nmFAFljPZTwJYxsLZPjtI3jrrEVGaA/WjSaF74rqC0hr73i7W1tjRMRILOm4xtp3z
ch6IX2qmIazHxg4/q+FJ+qp3Y0UeVakvZnYKjiwCh8f7JWAkPznUHwlD5Li0e8+5TlOsAghjwWpJ
PnVL6qAEbydRkyqy6wRJ1q9C879icnB1d81cUZAJE6q/c8I/rwTFfp8wJzx/WK9hRSSdTFoLUFCx
dxIB3JneeGmsGbEDFBRivAJsPMN6M26QrsZJA4gQ4xDueF5MuQwVlmpdSuRncodfnLgD1ohmWAeS
EfUl9JgUi8gTTARQqDQ9cy+Hgro7HS0atJ6JATjo9JJQw2tsY/CJULyYAb4pNWicLXULCG3AeScB
L98+VqG/4023eQBNsj1NP3Qzxqe3kIbPFPw2MYk7jurP4fAn3bBPh9Sgmv3fvFKNYbH2TdbqBP7y
3q9af6cX7qTc1B35gwPwggXg2zVVlaHJUUVB+jMgcVO/tKbH1ZjHesrrpOw6QXggQ1E9Wtslm2zF
tW5+fT8zvO2t/oYSqV4MswWS5XnMqObgLf90/7FqrBLa0ytaiB7wijvumXc1KVIvzSusXm/hN6Wd
/WiRfEyGjjKwBBevZ++xMudPZV7A4Ixi9iDCB/s+XjkDV1GWlV4mXjioOsv+kz4pu2JHUzhxwnwU
bF5Bmx1Ws88SKtuh7vaYsJOOXVrtqYFYIy57AAw1lHKSXQmRAXxeKFdRx2LyETQFhfXioxjNepLo
9pVtUWdy6UucHKyIaivGWqfOGvMLP5EBsM3lyoyODZQeV9EWfKPnTVQ6msvtBGXcd27i+U2Kfdwq
+r7nSb62tyZN8OblnxFfZoGvgZIEEf1GePfAPEdZfunghndavYGsN/8XELars6r29VRk1tYT3783
LiffYjM9Q6U2mVMTwoVcDQaESarCswmLmBUmzePP1qQaY/8FcK9Jj2zmEfFvjUXs6R3nh4fl2BwG
JwFnVOpMKWO/bTtqJHO8fAjepbE9YivEleSx0TW39IqFbrUjDcTKGicpBNU77k0C5Gdee+wEzrx6
A+TzKbk8FnusdnfBnruzupTIuV8KnKFxBJ19zqNjMKgFDyiK3SwQoZQ3JXSyIzWnVON6tybi20YX
ZUmhEvzF25FNKVUEh+Sol1ktcJxeCIUFbNCBwlfeMg9+MDU2jkg2QXoPp3k2xI3W5gKsriJBQV0b
bBfT6xajzJx3I5++UryGQcSo32+w40u3pLCeYUIJvw00OlqL4RRU1wRHD9j+vfbEGvW87ztmyY0W
7jSAtyQE1hXE/wnDB7jf72m35rMNn8Cuk4YvsOKg6BX7mWVBnYtnKXEzzA1TI90zh/NPzt2PMhr1
0cyCTpEFzUUwFZpHMlCh8c7otc7x2reZP9heBp+qtcI7cZALOKbcA5I6qJ1gtZLGaoWAv59zFtNx
nKdS+w+qI6x09L4Dfcu64Cb0Hg/cc0i1X0SSt+9Q8QBuTzH/0wWKOQIC8DIO/a1C3Mk7XnmJZthn
GuDeg223Yk1Ysq5G0mf8oUvtJrvLnQlec0WCHpOHaYiv49VY44KO+5AlaEgQ0gvF8aumwC6WjgC2
IFLH3Ym43OL9aQN7hkG3ZGHMbpt8wCJfF1xCLSTLTegzaeYEvQqLck5EpiRrbvywFm218Srq7Cs8
hc88eZzmffiMfjntEIFYKzQeOXkVczP8muD6HoMvIdVcMHSoZrE/6ssFQo08o29jyQmlyBjuwveY
swM66MW5K6o34xzaiQclNiXUTBVvtKlDL1xdY71/RXrmmOJgxU2bXYtnT1/Tgg8msRTG+47UrfJO
XGaMwB1/XpkSB5VxztSfo2PIYUO+phPnYYgpPj5ACe6y9RDILq1siMEOHYq8YqABioHu8KuBuBUO
NYYMSgFhoK5Vj7CRPNMfdszHyJ9KlAogjX3bN4rccauQBOS67OmfwCMFwROn1dOotiEswbZA+tE6
BYXQxVS1rhMdZdAwIvA50UjjQTR4sEJTg48UXcOaoCW7A3doez1YEyYYtrzGv9C+S9M/ex+iH2E/
RQo4XHcj/zdACjBg4wNXbwNmBQGyz0vnRPYy1gR4nF5tVfhi1s0ptBRXfoLL0uNcDGW1CnL19Jwn
tN4nOLaGER+hC1lB+M1aSWiEM9N8ZdTpEddav5N8iYZLDdbpLww1kxQH2OLuXnAa9TCQ5xPsTUAa
cDUGatUQyW06d8Sgw6HY8EG3Q+uDizuER8vvVk4P3HikFJGBlzSABnSCTdNF52X3mHrajInNl51M
7JrfR6EQKVeYK12Nn16wzpKLjcVhhIBzlE0tog2j7Kdzd49dicxlRKg9zMtn1U5osPIHoOO9YX3+
je9Jue1leMmbTbX/JNPU9Ld5F7UaJz+p5G9eIW25cuQNa+pRY78LH5evZdeeNbfua0sHW6eNWyfh
94KukdXjD2PVwHap9drNVaEWpynC+/omS6VRwrS4wKou/KEa8xjvfUjdqHYKfoDmjrNz0nHuw2Y4
jR21RCyW1xOjft5fTmoBsWIBBiaa3tNhSfwIKdctZ4AUTZ5mR9xZrvlcg8D1xzr92Seh/d5sveMc
WpVL+3S6M3fcC4dbNqxpMpIMHfalIn404JZBNsPfAGidSba04uRxUdJLX120/N5p8THzdDomXn9H
qdUjlpWlIdUoiaVsDTFy9cz1ShHKPyBbgQUKISEFrR5M7lyHq7caok4tqH9k3wDuxS9Qu9zEJCEK
fS/Zl3QxpsMh6c37JohsyUPyMIHVGuI9jfkbTwtufYC4aCYjS/RhkITdYVnk4/1yWC6z/NMaIOqR
j3HKrayZt1Bdk+Zk3qzxUUa/Y1Q93fwnPk/hI0i7UHcdbObm+jDv2BeGW6pqat11opbB2d0+GdOd
udupQzEzitFaXA8EiQ5aRn0bEDhsb0Nb8TRaFCDcHKEEUc7BRB7FSgBaE5V46mY9R2bFE/ylYtdp
yuLWkP/69aGF/PxoeJjxXdCnbzlEOoVTSrzWpzcdOp/u0+n8dxcp2ByENvlSxcVFNT4vHxj4OCAr
nXkoaPUbC3BwuO+koohJ9K6z3oWt72ccE1LiZj8Bj6cOCRm66MtFya5nQyW27PS12mfSqiuUkX5a
3umApcBXi8MLyxyiF+lxCoSpdXNwszLVJEoc7t3PvpcRWvZ1mODXZ3Q8N33rekw4WvjJIT3dm2AZ
uAFtA17Ic9nEQ6MP2b6aWT0DI+f+rjbHA+Z0KOkk06wGVZ7g/YLlBnotnj7d0JiC3wWtwXToaYLq
pG1gC82YNWFu+Lx/AzA8hfPnKOEyLg/Q4v7oKpI1SwKSQzPZko4w4IbjYK2hyVj4RC13ibfxnOfJ
/aWGc5kSH2GDC697oq6lMKtrAYFyX0nEv/dudBlOP4gRwYUgK/bnhHRQ5+C8Z2Tyv9x1Kc5JGVI0
nzkqVLFIIVSjpKlWWUXeFbjYXCzWMfLOgzuv+yjJ5aTh3JOzsezupRKdRSw1FQg1iBkq32l24EfX
3yU22KHOw/3CHu2eMsAEN0xvWTPpBU1FRlzExz5glDMufxy5q8Syv343NhDjWoELiCoCYaTso/Fz
zM7e7m1h9PCpzEJ2LlRJtfn2P2OEijtMtrVmlvR1SGYEpt//ubsOP03WZAw3DSxWqNwlNSGXl4H1
7NikLZwzHeIJx+kluP09RJPdPWQj+Opfhi5GFKkyV3tmw8eWWuA6A3J4G0DKxeJ+v6h/l7eJYmZq
Mvb/pRWBTyWLTvluDE+ojhV/9hnS3oxcOCUIJ4TMnZOldQm+pFYo24hct8sAxt+maofAIFLPNITD
LusziHB9jsq/lnEN3vMui1rZkmMZobd+
`pragma protect end_protected
