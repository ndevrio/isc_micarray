// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H&W)V^1,KBSZN6_6_7BL,+T%D=UG!\K2F5";/J1.Y+W5@P:AAZHIP;@  
HP/]Z?TK9BX>[)ZI6?NX1/K\G8E'@ZIT4(V<W"5AVZ (B6WG?$V@]W   
H&^F*PLM'W,)^O:+! H0BP%9?[,R?6XPR,RA/)'7?1I;]V*ABRJ4Z2   
H_FD!:0AS_ <=+)NWE#UDLHE0V]6GV9(@A#A!U&MZG;%:6=ZLHN5M\0  
H+TV%6+A/!<J<1DRGY;N2X++?.M10R/]-5U*T<?VWP%%Y."Q![8KEB@  
`pragma protect encoding=(enctype="uuencode",bytes=1312        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@2PGT]O0#^L %ISS59LC*7N_2X)BKECX?Z*8\?N/)W[  
@(/XJ86:KYOUGRO#BN9_"G6*76#F,K*(Z1$ Q"[S(?28 
@Y#R <(#UK;YOY# 8W-UV^P__;S(P:H0^ENV%D@)<:$@ 
@B@R[:(P9&BGYS80(&"-8W/%RUGD82P+-B%4*AS;]ML< 
@ZU2F)VUSM&&]M,>5#/CEZ/('-U/\;$[<: S:?6$0EC, 
@]'\WP>(6+?&.\V&\^?3:)3HQN*:Q%TW319]<-M &V3$ 
@%[7D8XSMSE%Y(Q7V<T^JFZ-D:'E$4E@G2R(:@(>U-/@ 
@W/D;$PI?L='&+.ABW< >?@Q@6U4^DR$&QEHF3W.(E@X 
@M<R 1CGK,K=[X=Y?O#W0-O<G.!,*:'Q8;*3IAVP<+0$ 
@'U2C06L?"Z6VVBGT9; <G"8H4!;J1V0/YDE'E*Q=^CX 
@J7962&WV2^>(K/PG=GHJ_BH7LU[U#!E]^> ""00<\\< 
@EYUGL=&7F53J/&\Y*:X+^[$N%<J+XN"_H6!Q+O]W0"8 
@W:.:294"#[_)KB?6=2_[IR3TWW2SU/&L&<NOW,@1CZ  
@C4I_JV47+Y^PCPA0P1R"I>V.WZY^1M9!?I(^@YM%C-( 
@2A.-G]+I6O8:,X#;N -:;N4HIG'S6ZQ]<W2KB]&7V2@ 
@1ATU2\Q;&ZK]&FD#203AH2B9=#NLILO6IQ9+$S0:%;T 
@QC* 3N2CLD&6/[\Y"'[".VB]XB@:W_5TTDR" WMM\5L 
@$9C)&C\Z61H^]AZ:XC>U&L!HU8=7Q:6;F?"#UCL ?G$ 
@17([#Z!XB^L?%U-0'EM4M L,5?X<VF;&;C^3[_X%>,T 
@>P4.K9C,;1[FY6BG9?:"A39NP*9:1IC@"^+5/1?M.B0 
@.]7!D8RO7W5.S+NM&%/.Z.L^,M"O:&E?$!M75C^R\4P 
@N@.?;WX,/P0AJ24?DID:[[J1*7_1<Q)]2D9/PXA#W9@ 
@AK".1:]D"YJ_9E$7->'ER7?PA/SL1NS-'\ I-1$4GXD 
@766>(0P=(N705U[TZ4=W_*.IVLVK?IQ/6G$!2A#6;=T 
@L[GC>=56O0&E'G]QU"0]84*@!0==IO"4D;O!.^DEF^8 
@Y.\<3(VJN;(!?(04]K1&X<#!E.U*7S6WII2LF!-T[?H 
@)"\N$9TLZ5KR]F"][J,'HTEDCR?C,+;LGNT8C;H=*]X 
@?9JM;:09:)\H1V[@ RAW@]2=D7T]&*"3[)<F&U,<H3H 
@Y.'/+YNY4"O4A>Y%V)C7.5);YW89(LY?M4.9:C8)/#  
@HW[XA]@\;! :D(7FLX,?B"A1^VSN#VE8)F'?U.5VB2D 
@.;->O7OM\#Q\K,83QN@LZ.7UR%ZTC._/5'M0XF$:954 
@&@L2/5#+.$5-G(QS>O/D&[)K]K<B]NDRS2>DQ86B(%T 
@FZ:.LE[Q,;6)+^XQ9IDWC*N'^=56 !:X,59M/?4!>UX 
@W/9^=$XKC*##04-3TF;..EAA@!TVQ%;<BI3K:I0L^X@ 
@#X%W]'!O^-L.ZC2T7ILZG1GFQ[/R+X#WFT/9&UC.(<$ 
@IO.?A@<:@[_N0Y&72N0:5T"O3^;(_>)-,OMA.I%:]$4 
@!7.H2,G5L!1/9=#-DF8S14E#M^Z+TNCH[!YI:AIP5C$ 
@U;WA#I95QCTH"9+/?ESEM6>G9^LBI(O)_PP59 =QT#\ 
@X,*MFGBW>N9MHWNQ*0&P?LD'IT>/#X^*-23 0K*%2I  
@(/;(7?C>LHOE2&ML;(T__Z4<^19"5I\;"S*#UV6[((D 
0?F2*O[EE7@GT7U16)]II@   
0BO;NEM'7SP<Y(&Y>\T$5A0  
`pragma protect end_protected
