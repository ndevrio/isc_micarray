-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
UbK59Wi7iUlFSHkCBDdZUa1j2yg6UY0fLJ5JBGhjtSxxGFeOWjZCC1zdlgF6N4Pu4Ykcswygg9F4
0IDEzND2lc6dKixak/z5EPISJE0tRz6/aQFGT3i9bWKWtBNebWz68F2dic/AMUHy+IijTA4P66XR
2SaNKNTOV5SK6tMYqvHyEn+JCPuSwYPbNq0xDcEmhizCUpdsoZGQWXG/x4uMWs/D2TGo24lNAH4l
nm/cjH8MS1g7GYT9qnw4etSC6d2g5u6y6en1gYiWUARdRCN9Wa8ls8zQNpwqd8l3r+GUlslRxumG
JXFpXgqEvyTmVt8ycNVUtXaTHAArYrPOptVlhw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3680)
`protect data_block
anE7TMlO1T7jkgFkanXlgbr0VWMTcEUq25Oy5EuCMmBBBVULQc+mLGunIGAT6bymV8FFxbebcZRI
sf3w361g3PQ+WGW1rH3BMP05a+ZA0MPo4qbchBJ9wdIyvIqVK0kH8q0Q+6CTki1/j9ebB9ETRp6x
LuzSjYnZE6TNzB/N4JWsIMx1A0oqpyL033p2ijyPMoaHxHByVg0DUei5WGpKSjhcQ5zmQESgAeZI
jTDIPAFHJjNxiSbOVEm0C9kaVn/BHcaKOhLZ4qKXLHTjTcorXfFb9vB4JTvD8L8axyRyJFIAVg6P
I+qOnk4ZwBWkbI+eyNNd8pN3H6mVRV/Ko1bPFhp3Di++9HKhv5xBzvs96IkeaVwO/zJIP0wogQiX
tsev1D6RCXO5++uyZ+V89hLh8IXS3Olp6saNXSSJU6eDJr/W+kMIvzznpnvHl7yxJqnDoqQC9N4D
ss932GQAleKtntB6raBLK01Gb2nQLnHUjchecngop+O8S7+MASXPZyaFw+MXPArxFxqU+IrpyKRH
D8mOanVKivUeP89iWncQJx5l8riHArKUiIPRB5J6JB1M/xrlCzuPZbqUNTSfr5SEKshi/ZAkV5d3
A/wV5A2ozih+8YjzVIzsICAHoY+vdd53iyOEZojj/hPNKQd1SutW0HxuwNBrxkx0s76QgSaguQWb
uBLVB6hwpXpUEIKv4kEYSvyFTSbs0/+0AXj4PwdBk+QUM4y0cKK7G075//IgKSy0yMq/jUjcY0Zh
XeBGrQFLK8uGg6X6XimgWlBRMy1GkH3R/tDZoiFyUxCNBMtGv16EGQlpBa8KiOYRpp+L0cH81D95
angQGzfbOZU6cFcRioX224C1wByXhUuiHQqKdCcXzM9GpPsLoXgs2Sfoy0AtXO2A+iyCjlESVdB+
8uY70v9YD9RzoBA+MlU2COkdE2HUTKSZz/h2+iU22G0kR8eANo8wJzpaKXba9pqyxAM3gDlZp0dF
Xz4Xp98VbkXAN0ksmNlf0VJcjqLIbDvt/k+SfBcqm+eZCDEBMddQ94qNDNaAzzjFx5/4foH4WVJ9
0b8Gg52Y6Fx7WXOjMYDQWu+CAgksIdUle9J7jKTW/sQFRtjltPrzR2u9sYLOn4rQCQXRHIFwMLH/
toncr/6ePPcY/h9F6gPeTCTZR0ahCFzV/i1/PKe03BYDeYgIvF7hDhPhaKjQ5jPi7kGmcga62Tsx
aSguKv4CAEYOrGf0+Lffco4W6/586cU9pYi3t1TrIjudeXqXWsZ6C+d8BbBagRyMQE0R2I41Zkwl
NO8BrWdF1ziE4Odk5oE1evS5XWe+XLyAStuGAiGg3txVkQEsRLHj6IdCJs/C8Tlr5oZpCNL28sig
1hVmxMnUWAcP4KAFxBaLkAMXzKGpOpEkUZKS8IIhlVvxdo1LE529rBwzAKNeuyIcmcJCbQHljSfM
8ojnfF8M32y/CAwwNuv14wg6MgFneK1rVf8juH5bo7qrSK3Lw2llnIhPdWd1F29+V6UJH3H38S0G
v1IWZTlLMWR69nGL5Xd66Tdbsnlys53hwnWHhHe8YTNERVbwqovfRzDwBn9EgPztbOQD+lcOw2cZ
vZubgFvyXNiQYKSQtlMm8rFAZ+GE7tPBYQAQk6UdkBmnMRyjxwKDcEbWyLpjFWHfAD1nxKPrbj5f
S2iWODN0OBLC26QCxMKTNnUpXsZ43Q7SM0ayXtsX5m4sWk8warV0Rfqz+e6ui29nPpo6GAR2chJU
LvwipeiclA3v9kCelX/WopTiKrlEHf0eRkXtj8xtqJGgcv7Q3B4C4U+10vYwOXsAqDHWylaoN/zz
li1msumHEO04WE4YHKryZnwuxJHj5zt+sLvMS6n+8/U10c+mi/g4Pt/e+TuXYYGNuC8nEwsE58KB
CCRvN1BkG6nJuyv17bB/Enod9AJ16sPbhBIZxsQwWpctY0iyLzdUdejNg0DG92aQl/ZudydlaUBr
GumpFef4SNTRJxINp1g1Rl7asgC8CrC8oKseGC1LwLWwCDxjUrF3CDMy7jsadDR9XkGu2zDyqDJu
w4QX0DZy1MsW5OFEu7TfkE+DuCLxm8hFoy5ORmS70/8lghPoU0oQqfK4C92KtTao9pPkaPYQLuIZ
YBHXgyMWRaJQbWTTkvxTQ2upPsx1POEI7Mv7aqe8WqhLMHYq0SPGasg6OQdw+KbwzWGIWnrYTV7g
+XYj00YFgYszoY8TzrQJH3waBevft64BafuLfoz12tBC3x4cPSLxYU9hnet9MuPjOUqO70ZZKiXz
LuZgTQ9mUqEhLYXUfknMEjko2jPzXSpZkuRVEo8I/yh1ei4fGHjFzT6WFN90muzQ8jAcJ5yLD0w3
YrQSIFm/52+xSllBA1z+aVlu7tE5OWv+3y1yBDWBB0MYfq/A+XkV1hyca1kAGcWKwLlqgALw2UBa
rKvVNrqhm5LMEIrfv6p9QJUAS3y2uhsBJd2/aPJzTs5xyiAXqC+cNMRdB8kby6PWZ2LTB4p8nd8s
g1WcbV05M/bLV/yz2xsZHBYkPgjS+i1es4NaN46nbjmtMNo7Hy2tGHBHhaVssfScwM+GceZbB7Ne
9h0mt6aHlAkCNpEOy+b+BnTxYH6XnjKex8eqooehPKc32bZ4N5ond8Pmfscxtry5RFevDjfvjl4W
LZweFAUxXooDp8AZaIFiRj6xicHAgx9wN9QlbBmflM7xHiwQiCWU/6Ftre3ZqGdW9GUykZrdnQI+
9aMcfulv7MNM4a5cp7oyaZMZVw9jKNTYLXWyy09oUBUoKqzAhUjDG7ZeK+GUXrkXwgLL5FtoiSuQ
xfeWjIswjQivju1OboN41q6/0qaQIjthO6lqd1yvLOq2CRbRblIYbaM3rKqYUoLKHfqAAwYk5O/3
SqmXTezx5JXAm2cbWZuja/Em5cKycPZkljNrsefl1DJHHE/2VyRkzytMtCH+bnn1wIuvwy/7EhYU
hjXcSKDNxt7lARdoYX32DeS4dfsfGgJWMDgGAOZENX0TvAvNG7NZwNu8n3z1RAFXMCc7bYBdkGBJ
wGIxWCkqPK0bTqZRbh12biD1hB9DUEUDJ/Q+uAVIBtRIB5SiyzfGo4jkNuNdlgLnp6n0o8FHsby7
Qzl8gKkj7ZSLAp1pKluOW6Kqp9Wn9SP+cm5HBZOe/g/0jsEtRM9R//DRMVql+ExA/BFNSXKTfgV6
8gk6iTAUwJhXNX8JDhBPOk+CnCO0NlUGGvHz8pljNmmpcIm1AfLvYL9N5Kh7ben6Qy/8IHwWU0N6
JQXUf9Pmyeeas+KxcVrl99Im5Dv0bqSFHNablxOzV1deaA7ae803tlBS0zZe3pgfMyJOXMZw9CvZ
rNvysmPpHwf0MAaKYZ0E0ekRGdQD//B2jTg3QY3HY4H0mXuh7OUNLvndqVBtGvJwrCwfSEdqr0NM
IwbAg2sy9/pEb/C87yGyBnKSP8cBral2hRWZzuUJs1WsrkT92zXadw803OujybPtMvAH0JvJPj+4
69dZG17woHUl4swZuQYAMbft4ta3yrswZTjqxpkIDphmffX2SmkgyxoBRPQ+e5+ND7VrKTQyNm8s
pjMtP4aI7Mv+EavN3XmYWcXhF9HILHD6tICrOf/ukz1nIY8UfzvX83plOfQnnlJS5STBYZ2NUej1
HzGOci0+VpfAbXxy8T3g2pj7qp0jE3ffvpna8+RnjX8BTRf9iETa6hPnxKD986CUZfVRk/MBHuqL
pjXebCPtwesWZazUPHqenpuoBKOaT6zgugMQViYq3wS0sNWzkNe7kWCh65Lxazt1TpHVqrrRWB/U
+YFKGcpDE9GZsFBn89yhn9AJ34wzAZllUwmAKwD42hHpl7A3jtp3PCwBczE2nBK/iD/57jBBX0aZ
ZnKeWnZ1S6cYkJ7P1iVas1fSJB+ByTvRBZ8bc8Q9JkGSGDtdbh5YCnjaAw19SsqefAf5+GGZEe4M
bVPry3t4V5rmv2kCTzMdhPRgDSlCxjCaRxQSdBhFn4+p0AlL5qjR6xysG27ea7j25HNdGQ5daGGX
EOR87RhpSMnQ8+UjR1yIxkp5X3hzRfh3yhhP9nEv4WiRBfg1iaXeH5A2kM0omo6Nk5/lrrUeU25s
9j3DzLWcZ2blwF6ARRsPMKyvfNUap4eIklWD6T37qAZyPYlBviMCp2tDEzzxTYeos1/ysQZ/qvaU
LXRGtS7msy5m5V7lNFCRgK0Gv/DTg/QWxzr+t9kYgBup93yyIwy8pJ2DP6stEA4IhgvOVCb+xsBk
Q29oCfFMHzyd2IjEXpIktrA+sB5KlV6harwKJfYZPepbOPoSYz8OvOOL2on1jWRK6bqRWUi6c8Wf
12NBBPvtvg1lQscWax4NBJV5I5DjDH5zOrelpFUTIpK0hdTad1LA1JkEmUXirP64tKWrf2FG0tp6
tWm1932ISn0xsgznUBpRsLH5omOdhD0k0RVyuKGv98sUhBDWR3J78AKKIbRT82gtCIRjHsrwmWDH
yh9Gjb/osqSbI+DYHDJp4sWa2PZnDqOQ1PknuQd+GXjiucCCJkSRzNYZJKKxgc8D95soQJ1WfLKk
R0GT8VzTG5t+3benLY5Eab785xI07IVWvyR7LTNcz1YPOFt+7ab5MJX0LW3wtBXWuMny828Wqcq/
OmqZd0ZPbgahUP3O6gjja6Tc229vhcu2c2l+7Q6oqsgTZ0WJKxUi37YsfUzJHbZzMFejtSXOJa93
7MHx0nuepf9F9EwQf0yArJyH7UUIuJU11QJ3N0MCQlG1C6pPknM1krctq0Lqo8IubKu2T1+OGE9O
+eEibewVObj5vFTEHQth7+VnQWpxDxQHHu3kjNbMPiIAPY2opMXgM/to1YrDdhdDbZGSf6Jsn8m+
EgYPw+08CLxBDgzVmpOR4irBy3SKY5tw8Jg52UpEcnk=
`protect end_protected
