// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ry1TCu5mDHrktey97nvF2cOnozIDpYiI3nuHnZ+5vuAvr/mLe3WjZ1EwWGqvWS+SVCPWR4e4vdlc
w3jIdUuf4soXvTfD6wHmd69C6450PwhAjtBdHsXA8VNXxGrXQbIbmHj+XbSK1PI34AhQA44lni9x
u0/Qdvhn3F38N1OcUQ3t8GyADrMrNOdxYYfBgw1KHzZXLwTnsTFQ7QHToBd8VNTKMDv574WSkf53
6gmCWXNeOV66MpKMRe0ApG2aM3c2dobtiWG2/9peRmOBbambh4sIDWAGfqeLf+PJP7rCtVpAYbF5
5/nA3EnTJjXttVvgJ6cmOtbV5LJzu6WyF9BXkw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 22144)
wKKxFf3d/XM9iyF01PH3Tk0hGhtRQ5vDaMK9mh15+r/UytLH3muMtDI1J9Q5QnJKlGffWWtTMjOr
ElGVhFiYIqsXgw5D+pCw1zj+BIHVtmsf87QFKMUk+OlPdA5thPsMuPQ8qI5KXa3QOU98Znx88Fhm
Xh1z5Dtl+MRfqp82LUph94Hlu+z0MpyAOs+ivvRgXQEllek4sYqhe6+CIyhgS0N2MOd0Vadl3Emz
DxIazVELcBGhp26SoCpO3BkSKSEkQq/kR5DxbImDWRvLkx9PfVFXu6pjGJLzIh9hdbPzIUY+Yn4r
oOFLB86Zo4H3XI14hdf4ctmvdplLszUNSBolrBf4k1AVYOnC59IpFcVUGhcFwE77qn3lhY8oTeUh
tie6GYhWInv/sGF5v25zPHCVtK66UDku7GAg5TPvH9CkI8KLn2gT3g8n4hTkzllfyzrwY+6Oj161
ZElDzhaiI+ptt44qYZ6nFfGlDo0RbTl0XN06FtsgilMK8pKJTqipva28UBCTjsx52QZcVfeljpEb
rQaEHjMh5i9TzXK+AzgPUsQpYgbJ5ChtM0FuBbawosXbdaiA2MNB2Bfw4q+q8lyQ/vrWUzrP6/5+
2KkjdGy7vw7Av0AQz9GAtqnuAEBSuTH9EEAF+EsgKvmwwNI4y1P+tjD/Vux5ohD1ZCTZxdqVe1xO
zldwEmzNs5xYkHfz13vKhn8Hui1tn2f9JY7/ICoQrwuFmXftzqHR/+05upxEK5adkmTymz42mpTP
CINaO48T1UJMWgI3dt/wCSzfEJ1zq19guOf524QqVHXpkQCIw6pMb7h5S0hxRQ+kv08dHDgI/ySC
4m7oUad7cnlKw+1izVuX7Pf0t58e8Xwy289u2uPu3+Pc3Skk3z+peWKstGNIR+RlA57UG58O5gcz
ZL6kyzzRI17yBJGl6DK5WTHK2To9bpTL3KxvFYyen4h06vYNfIlGxc3HXaCKF89EHIzCs400zuD4
ZVpwMerNsrOE8yWS7iccMrtJZYQDebb8JTzNDK0EW5C/aJQ0H3ylrAPOr1grC2XE8BPapu1k/LX/
0ORWvf6hZOg4UBjPk8wJQmjnk5Rc4+/56vMEHUDcQfnyDDDTPxJUcv+eFRyI6BMfyFL7/BcvvzVk
VHo19k6W2Ikn5DDeWsfFp3L+avSO4Rq4VLYuMRpbFuNh2DJW3bXjhU3nA2ZvA3ufiJ+/LsyavyYF
kw84V62MBrmH0MX6r+VqTI9Mo27rhVbHuwSqs/5qCvdxPFXxNAmIZ3wnI2o9IICVJ+PpFORCJrxA
SG8oUR8BIy7BkimPHty9aMtYLjWbsFBsl/IPLo6iANGS7vtrzmbbTDP8BianLSxrynpO6MCFjiMh
CuX2WJcvGqIGaFIh5gSJhde74bnXK01T4sOKrkOjKQML24QBJFrGd1E4xjSo7MYp0xMO7JG/m5EY
e1RJIvbfAtkIZFzYCk7F0edQdmkJy//GxiONL8+ipJ2MvFiLWxkUTIuptYSvRDigtTCDoA2WKL1B
I+y2H8etYcRVfqIHH/kl0mJZz0vmcV1pA9YPzYGoiS3s/tnSbEntn71Fw4UH0Gw7VNgZy9GwZ2MM
BssajovMBrbdbZicXFbIFbgqlA/uOlWSuLlhks02rRMOKZ5SwQC/aPZ0V1jiZg3z9xHASijU4N6S
AUkWPm5Zcl2QJXehj8cdBDV7C/r6KIVGafb3/4BQbMouDpvnurWgLOXVtmD62YJRWFA4QTGfNPrj
gHaBX2u43JAXvzZ4EkcPT3AoJINxiFt85fr3ZJGlSxX96OXzdXS5/hxL9695vxD0uJgcBWiffK/B
9xIqUdAyM2Gfcg2IDd9caji28dAza6iOo1mwa6sKSih5qLERifMyXX0JL0f4zWFb23Svq1XicRlb
JJJjmKFr1nc1auC1JwhUSXdgJIhaz+hDEeeZOxEzWFlTB9hn48UJlNeGUZOUwbsVxkVGQbZyF+FG
YFcGV1VgUlm+qMIwguw7e697XWMahWsRynw75fIRty6DepEuwLSjNX3kLiG3QrkJj60WbTEgeTm3
jG2r3zJmyVjF05sE/JAgNDJMw4KFcrFWm6f3JETsuRN+CS+JlsZVjMKc+RfMMiELqCX+Bie6TFp2
YUlKHqtbT0/BiAEElY/BdKofeU4waThlYcWMX9hsN0XzTSKjSPxizNstf+vl8cPqv04v3/sFuXSR
FSWl4RVGK6CDcJ1vF1+QAtL4prhCSdGf18yRDD3PN6Oc9lsKbFK4Ju5J6nJ4VYchtBMZjq0jZJS4
+BP4LAc8e7baHCdMcdPhK0RdPGi73mVWgXcPzlOnYFwoWA9BV75lFf+9O5fosetnDK1pe3EMJYFa
RBZKaLhl8MlLdt+ARED0QCES/iuK3mVSKINrk+ulsLpRGR6wbrPD8vcNtwX2EsQDMNbLx19BnnDZ
qc/IM9kCNH/co9vMdJr0MpxU+y9FAfMGdzhYzADQNrMWPVhGj3K6rbduUUjQ/h+FYhJnCUuDilnu
qQ8416Gfd6gpj7k10TCu4lMOo+sO0cd9Q/zEI8G4aHstP5SnGOypp5Gg0duWZaoXZ8q1DwY/lDvC
Qd2cI3N1P9VNNsjDwVjw3aCHpOksxAocqkeV5u6IFlFAXKnSUvItOIBDN/TSTCJMDY2euYoAoWco
w3lpa1Lof34JuRRjK1NJ/fD/LrhOmzdDsy3fapkua82CUb93WWaf8/jZB7XCf5ZrVb3+gBcmGM1b
TgBB6/CI/nIt/5315HID0bi0GDdzdLB/bbHzUoL2zJwqaQnTY7ytC1YiPRjYsrGIhRsypaQUj80N
DWuCSFryVhtV7XVdQGtYzSVWccGLj62Svpu2p9EKWoQJy7uhBd7JlG6jnwSyKhoIoOg5X8xLQshv
YowGoFnUUG+P2C6By66slMZ8dEa2RwgDv+n1IXJXjCjMAsqlotIvhlV0w+TaLSj6+cz1dUsjLS/t
VL12QUACeehmG9ByJG09jrGP1lutrl09ZIYd9OpvIGAxKUpl1Pdoigas7JRxUnX7o148Plzk0vS5
G89JIg+QQYvmr+rPaz5Fuk20cgQdoHjvgUlbJzRqVpnLJtdPEzMDTPJzmtFkKcMXv0uS9U9eiR2H
fKE5goz0S3LrDBkr6ti3gzv1Mgvk2qHHnMfyLx0HFkJ4nyhxxxkLshlc+il/Q8fOyWzPEUV6bDHe
rnyvwYwgL4MLkSbLQPE3zisKNMb14mwuUfWpEJCoZjWvI39Yokx6IECs2nN+xWPqrxO46dMOi8ii
5m+uenNlIzU3fZvsTU6+9aKJiwGWtTdQ8VxcXIBgOYvk2EmTD/ubbcD6O9KLgGdVcy7qz0SUH81a
TYpwYZ+C3UKrshnCh4Ap3PBmAfwStdoEXtlmVz0zr6lEaVCNGoIsQ0B7N+smUVG03cggEvOd9LsP
F7mqlEuUiN4jT0ktdsZsiyo6DtLd0vdQoWcARqCHUx8NHOdZfnwb0MKnnphhbDV/VoX1MKbUwtVG
RUdAN2U67GY7oDgl5YDBMOeqTxF85KNuhxugAK1VdsG/jN6aLiRbaQLgLM4BLBScu18A4kss7Qlx
93qU0EDs/IuSezGDdoyJ+Zh62Kap45k7eVci3FihUojaA/dy9DW/OPavQG6iwxcA6esctcThMgMc
vJQ/Z9CVGgX8UB5XOpLBrZPyKtlF6B481uGrrEqy9xKAKJdIi3367VnJN1qp1TiD85hNWW+KiKj0
bqxqrGFT48v/Zx42dSZXl7eSEDOC3qb4Jt+CYrUPpGVtGcRvC2b4RdS4IViUFI8kp6CwwkFdB04M
6DR5E/M0WCJGWSWTTaZsyEUuo7NtZxivVTJKura1OYpzfLz4ABKyzdIQ7LCvPmxJMF3rnr+Ahkit
UGlFBtWRkpvvAiK99GcTfL6yIVVvqCw7SGyQ/Q+rpTYpOzu4c0jHqMlCGknn/HL8Wc9sdLLU9I38
Nmf/sIjRTExt/8xwhOuSmsrP1kCgBJHwFcL1WCCjKoGRFSDKF2z5KftrgQ65z+Er/4De5kk7/qLK
YsH2szIWq/ulmoKQ05y6eSX0QC4ypUF/Qd5eyWCeTmNVY8+xBWaAvlk/XlUr8lrt0KglS7721BW2
VgQKACwXLyMZmFDuGiE7XIe9XbNm2mdeNJ3Y/rjUVHN58znDzHWTVNx0BYxE0IYT9P7Lp/qKwBJY
qVnPhRf3Jg+guLrl6i3CiGkRi2L8rDhejLmuY5AsZirg/yAkIUuOQALQ8qOOeJoa3hD5PTiwdhTg
YyJEUs79opgresrpk6AKGwCWlpeKKuCrlme06aPOrQCZHASYlv5OUahbkjdbDzghnFE/VFiM4A9c
fI3o7JzlD3ju3mvtlw82M1oaXTby6rJS/gMUTYLWoiy2u5vL5PEQenEnk0Yolw3I3WoZgIN+ES4u
49+Rt3Q6GvIVTvCB+UWcuqT/Yjx1viOSLi5Z66m7fZIgU1AOIetbLP/9cRuSY9MG+vD5lAuXKBMp
FGGQYmoUGIgXKNorGyUVcnf/fi1HYKjquGr8+GPXxCzMN+Pc87n/6/c5H6SpFHwmtne8pmcHPpec
4QiJ7NBff5kteyTSGFUk48TtdnrCAOpDGwF6DUODwsi3oOSP+0InEO9sgww3jh0yZ7UH+1X0aRy7
bdeEBTa8lU3CnSJUHtZ6VYyhltrloP3JhxQVgFNx/TgM87MSmEhHSE1pGZHRB7ORecm1/DMvKvzv
fSzxKKLvYcFBM8094tGtegceB9RH5Bchxq8V34STOmr8zwSdcG5dCxYcsBWBFEdndvW5LK0vYOs3
P6c72+ADXZwKvq7GSPHnQnMolXpHX6fB4WJHEuswd9wPDqM22wVvaj5Swo5EOyLiUbRsc/XkRZd1
L2Aiobr1sUji1BY0DKfuhaOPk2/Nf8SzULHptbqW1M9dMIaVDFYmTIn4f5of8+pjr1PZldbvYMs2
FQIogpN6wrpX5jJIt14DCiUjYK9tbNw2Icdba3Pb5ubUIA6utFnp3p/hnA/PHjoDp6xCZyIfqLpv
ZKXex7Ndoj5Y3gQ7voIz50Oa56xp21mNKHUVN39cbA7SG4prVWqmxCCnS8lAhRsy2yjd02qIMLy+
YDb1cGG7KTrv//nCByVpwoCSTlG5kaQtmj6GOYzXgjEW5gN1qfPzD3f7huioiX957E8tTmM+Apb6
Otthbm1dWHGPEHL0LR0EAEK5NP+pIjdgj8WaSRE11/f/gXVm2txtWg7qmfwivFC3zc+X4bB7qlNq
AZc0iHe6voOe3sq/aO/xslgc6xELqX1I+m7fwERPE5NIeOEHSWIVw5hUywU+GjVGTH1TyKNf/5Kl
d3b5mv4Muft8U4HbDqgJdyLPu1FbMeqggUr3PNp83QUjlaR4YES/Fuxe7BzBSNls8edIBmz0kJFu
CDp1NJkamvr5in8DD5N9yts7qY54K9iQ7tVB1jUlXbQLkICO3Wj4JSw9n4NnsShetKZN1+9u5C5P
Iwc35S7XtQpaRmSd7xFUpbNRzxQSaW0d648MO4o0dLCjFkAWdJgQs3ftntPjXdjZgB8hASWjhteX
iIt9ER5lxdrT3Nt/7eRfzu6a/8eiA2KHr0cZamPuZjrbAWM5MnuJ8V066AbMYSZhIRsKJtLdzKkm
WyMDSuSLQqDhoT5XfGiHFSABkzt0sk0RXidG9zRNW+kOZINUa1QdafklwvAX321JkNxXCIZEMHT1
kFy25WoGfChUwM7/6OuUfVpmsAwLFHjf7TpPNKPoqHkQggthVwzxt/3oi1lVxGHznbZebeK/xUyY
yCuMPXreK72lTn8HLXWqN9tdukVMZyRtUbEmn6quT0B6imycl12/E1fJgJ3WSmcEASPnl17U3N9Z
+PbmEIAg0w6jmWrBWQCYZHZ5Ub5AWf1t+gpCK+p10kcaDOAm254lP89jnxq0HyN1dg1uLVG0X86n
vMvDUbvxRkPIG2HNMJUfXbFlRW96mnVFK7EL1EIqMPA8zPAZbIiVg9rIDPrV/S5SmiSkRNhbnyxF
Q0i2VPFxVCHRkrJQxfSWqglq2x66AmObZmLwxGR8vv4Mvx7zBCxTXeyG+sQraMbsfDPjxu5wTZ+G
Um4/W1PDXQtQaldZM5ksOgpQ2Y1bBgAtNevJlkMNOhNye/c+koyZLwg64cWtGjVVS4ghOqJevyU1
aZQEtve4w3M4QxQA+t7K+W6qGQA8emZwIFJ0Yv9UtUGV1plIFhXbRG9TXh1XR40r3pZBftlsu249
syXO4pO3/ZmyQ2YmsST/NHGi3wrUgfrVtKxRS5ZgbpWsWSX/fMZTkNAEwFTqBdWvN0zS2+RQZKCB
tQg0a+ry+LAJU7Shua6kbp94hvv27dabte8uQinfwvHlaIxlVUT0GeLbRroI1wHXcI2njQn5ZWdT
ZDSo5fqsgjpkeHqTmoCbje/XKhwQbNycz+VNhdTC3QxuLthX1S4DzHsf7yo/2cGPBLUK4V+0ygyR
maMSl5Al/r2CLMaWnSvMxtxjahbwW59YhGidZ614zLsM3xZDzjg/8HDX5TMs03W0BhcLqzYSNhod
HJ0+m0YXpZn+XZLi0NPSLNRZG5cTSo7yVsYXkeWask1IldVWKMHwB0U6574o6x1TbwMVb0+5BMB3
rJVoLmbPjCSIIKi7qlJjWtXAa3z+T1HrGFi7kcwJcZKLRE3ZUybDuTd47HKIkPorwZ64l+oSOdzE
OpVBaZPo832RTR4I5ubpTkUQ9spGcnkY87iRsWbwyJlyrgR8Q4C+giInNzGb4LT3sHNVBtOMqDHT
TnDQ9Ps1Al86ZUmprYFCU+WolyX7dpXtR+q+WDwuLXQh3jAOiIc1IQNE4ZtZmnNa1LjaXFPyuVJ3
05XXhDEBiannkZwHOZLRI1GXvTYS0IMkYu/tWl8sAbNyExU7Q0hm0daCjmN4miKzO2eTqpBZjdiF
S6LD4ZYNjLc0czb5EfnuriD+yv+FlwMn9FbSg/qj4WQzKNgh+5W3BeKCl6/tVMXnRM+RqG7vPPdS
YUEALL74zuRF7PtfVqMvMdvPPmvjApQsjQwd9w2Wppd//N8LCs5bTNQqiZHWVlDc75zK7JTeSpED
rZ2GeyGxLSbcxWo+3Flx4rjpqa7jbrUqvbtl9JHQa/svR0gSWiecGAQoI2IJV6u2EEpYyOd078z8
caQqmnyHeKK83uZvP01eVw4RTEhMEKYEwO0uPJWvCQVZI55mf5zDHyNvpp4Iu9TOvX7AsJJodWOa
LwEmRyBNh/sKkg29qGNUxVjTJsr/0SU3PU9d9eSsB+7kxJyeGiXM1snqcnBm0ts7C3GyyI7sXok3
dci3tDQ/kj2UGbgJ9tAkBnDKBiILyOq2mDVzwR+auWkPUJ1K2YQDmY0yxUojF2dGuItPUlPXcFoA
29LHzFHRBM996f6raTF3KTqv7EB+v8CT8SJ09CKDmaqtbiWCn90ibLoQ/k8qFKYmFKR/YbLpCNtK
OPsRksKjpqos+cr+/rwuGwP5VeZi+lDmR16o2zo9lmjSPkP0JG+EzaLYSlzYKINzSNYKbK1zzEhM
/FteZYVlP73hfOS+sAQgcKXzgoyh+5vSElRNCarr78zNjaL9ycI6N2zcwdoRIs7ltBNEoMvrUQD6
b0isbkKZ/P8gqFXfCBP+/YmHkZchMBfc0RFO4ap4Z+l8BtJjsHIJPUVP5bziVOxY7UXdZwXj6fv4
/ICgMTZ4cVcfa9dFGU66N5gQGK//E6Pd+PoX80EMQugHpz78bTvGPGq0bJKuPebHJIznC0hD+WR4
hlrtcDlnNLXJENWcjRUyaW6jgrvyYXO7fcqzrPRrXEtbkpZoHDG9K9M5nrBN+k4OOZoRdNTpJrQr
PrajeLQ+0unPL+8FtKkXO22jbwoKNaZeWUhOs059Tzgwr58xSWgqqRm2VnG+au0Su7hyUvUwUA0d
oKQ5RC7bkFZoA9xL1EAvBrDbQsElo+VVDyLp3japA/cYKnwycx3qeNfs9bRXxFE2BV+LquUZkr0+
6+rFWKMgcMgU59A39pSRr548xNzmtcvdJVz0CrSrZutkCAZXEzTbiy8pRKG25SGueKSRjkc+MM43
DJoKf476bOF/n3za6Qf1uYxRltNUXSq8cZeE3wdNX6hwXjp9johYWzfJesWqb/Awy9NvHU1mTZV0
rdvhYMnNjsoK3bFO131AQC9N1fSAM5fUtX/iAH1hQEkiVG+ozNIZq/P3t+GbUdsUadThSjIUixEY
HXubOoUqeCOVGwXmsKyQp4E19a+Mq5pOzPU5BztttWbiCw3flKB+9oGQ83959a50WU0xwlWaU2eF
QVrTsV2+MlC4SmzAa1+hL9198Ep67uPohNaMTssBoAnSeD01DMvsIdtxu9ri6INNreN4UCi+JaFe
83bQJxwGx/Ag7exK9gVbcWaSILwG03HKC56/x0Fc3f9pqv5n7MfnZOZE0WsnIh5Vb4JcM3oPeVHx
9ZsBNSMD5uZqDzv2FlQadbvLT2sthq8Kmit+PUNoNceQx0giC0jixmDmUfb65F4/vPWlkB9VVeFb
hFcHL2Hq5P0bA3cTgekImE+kZp3Whq5IdBSx0oU9e2gGd3pwYa/3ebWEoynyly0GLL3MHQccBpgf
tN9tO7xwAigtixNI+PNoHbz3ZlIrpTbQQDVbyKaDTcD+j7sQ5QYsnvTb61MHzx4hkUeoyfg0LsBC
qViFLQcDqvOUeQLccPaZy0BaouxA6jH0d8KfGENUH4j6yU4ScCfB4qlbghjj7KNoaysw7qKq02AU
0DDlAmmeQt59ki4VtEqmQEnlNJiQq+416X8xuxZShbA1Xchggrwpc39Wqe/u14fhziBUorufl7f+
poaBYwBKyVPfiBwTwvLSpfuqhqowhcLMg3t2mwZ2h6iiLJvm8duToM7DAn3ohljXqHAW1x58hUIf
5G3erUo70QfsygnnAOW+ukZs/9CB5vWzX9qPWqRYfiJ4zEbczCahvZCef+nGHpb35mV6XAGzdCXE
tuFQXNm7YhpzkWy3cF3xdGP3vYR5T7n+n99Deqeky3BCXKDiU8Aj+14RPFyEh3qNk4YqfYrqJQYs
IYiYcATCadnpZuPic9YyCF+A2V0TwxFkSkrv4cZ86KdwbSKyNrb/ofe78kFDRKRi7TTk59JvtLIU
vByEPeIEKDl2/NP3oZlKtiDkuIU9jblDYcmxHnBRaXhf9ZHsjffeDSGua0UO/ZfIwcSuZk6hnxcl
8oWo7o6ecZidADGQYl6E70w9EW3MfBjY7CDR9fqx1HSwfXYy9qXHqvZ14OuOIDABlzfegu6EUwVO
2/XKsJeEP33EhE91gzGQZlMzz7q5RaEwFIjNg116L1xuZsxx0skyFILf5f+o44DnFr9HNYSHA8QZ
AclCGTcJP8sK1fGoahUC1nUY2SV+bln88stL2WXGNyASWNBB0aSkNOzGCAHiDiiUN92nCTuxU+2A
S39Ia+58/o5nnK+nOIQZk505nWiVyhedBAiQZErgH7pEnl2VSnWSOw+x01bRouZ4y60qDPFyj6ez
UL/6KKx9ucbYvyNbsaO9Qp+sQn/qINMVdOeFTg43mUM0gVR15ily3HSleZ8/dmxb3cU7P2IhOCsh
XJDOgeS6ptD1XMcZzd4hBPKHRHzP7m7x8g3+0BWLhO/hosy1YORvMaQuKRFyz3z6DbnjQdduo+bl
KHoMmZhLmDyKAjLp/KCpatIxVYND/Rnll0gHjf9oswb15+XnANx7zq1a1j45HuuMIwu9LIMea//M
J9SZsaRvAVjDs4ZtC781cCu46jGBKasPt04Rybldq8E9gP9SezDHW6GBD6/bKyulxHfKK9K3z69m
vxmU6TC8wqgOaag/aYntCpmDbuuVgYscNJFPt4ncGfyoVNQlTsarxWJbfCP2MrFtESsBWxAzE3BQ
MeyJiPTOVdzrMfRKsUHIsQ4FL/IpavZZLvlCLVbhQHkS7tytR55+H0S5jphGUXlhLQDd4DWm3jEo
6GlYqOto00iHyINlcB8G3ZKxfXEtUd521Qug6ahFXqMh9xjRdDIIcOcO3g2nm+X5o1oMQyNquOQq
EiL4g++dL2mwECWpE719xMCsiE3xEdmfQg9bpyEl+SF7SIzmYw2GY6E3y+sUCg7fm3ghsMB2yoSF
Sf3MyzZDSM1ktRQ+eRvPP40tFGVZbL61/eOiDXN++z5hbDRnpTIqYToqPZP5IMSF7weQXZnvTvDj
IXrfehCAJ4Bqv3k5bXjQGe0VJHDHsUmPALUDTeX7dnGwvl/5i5mCXO28qof+A8zHaWhI/DuoMOjz
hGRFOVGcFbxMFY2HnJZfiYMWoEaDTcvXPFrij+MF/4ot6jL84DIBATufUliKRgiaQR0Jrcj2GB++
VPlxu0McZ5rglBb1P7sBo5M/+n73V5xIe9Mr98RqKsNSPXZmxL/22OnfkLfxFkMGzYCWQU5HXgBQ
V1dxrH/F6FpP9s6/1HLWMuS8BizNwboWC1J425p3xRVrDLFp4lG3KRKEWsOa47Xlv+rMVQLe+sjt
GA4Uo26NwfIUT6R1R3ZmsVm0Mc+V1DNuxJQQMzGlgDr2aVJr2P3LacqclQVZGL13wRt0UZ7ifKnn
2e39DmLR4ZaE0HhOvgoGlz2Wtj5gcVvsj36AlwvjOZtv3hiphqnP363jHIwJd7f9Ol4mw5HkSgAq
Ns3t7rhTwwsvCf2ugDCrXUOMjtpwsLAvpxZG4eabE54X+aDHeuZ4j8xc4rjwetVaiw3lcuk9kbHw
vnApvCp/TWcReqLw7w+vguWZ6WxAG24WyrysOfd3icPt6MjvOtBNSzsWHkIqXKgRBg0u8ST9BMRK
1DDVZxUfgmPnih17+BKvnLeWokWLJQuOu1F0LW+sOl/+2zjlyfbcO2aEsdcahTFDGQntV+Fj+cf7
hvxCkgM+OSkh0853uMXECvRrxj95lL7ilRnOSufSq4Awir1ChUy5OLX1fyeAAL54IvCCjfptts4T
tYxF3Q+tdEJUt0Id4d8IJ1y1PPNxh6QXD4HBfwrv/RMAoAU1B/KS9Pb4JuTU5ttGky8Wzwrl+Yug
79u6htV/c9sUNamNnVgEnXrMb9b9D2eEmHo5uOqq5ud9ksSKNs+/E/m+mbP29Uf9dIE9ytoGgGup
JsVIv68FBhcqxpqKmqdfBkpZcOaWHQwanzpb9yNX7r7NUggRtrABaZV24ulEsJbNpCmhnh58k4sN
g8/JPfawfoUZyt6xnfcC+PcdjpWpSOmxa5nUcUhV04iHe57Xe3Xs7gQsDsHy9TGheUei4sZNMUSl
7hT/GJ2Q1BO8fPI8obOCnah7MRfnaZkzzqGo2Ru6+XsaHOtlkk/qomx9wL+csN6Szud3xJp9HIOq
P93sqtHn9/AVd11ZJf+Ex6w+gGRnfb/r5WXXj7B/DGmy0zuWQ+080NZhLQwbnmPZ9S84FKkmxFN7
8JPj75zXpjTv6weuoxvJCFkEgU9BqQGpEjDvgjvJjh36eP8JzSd7DzKAnKuKgKkZ3f4QVlKJL0a1
k3kNYje0ley/wC2kZjeJGKkc1DHr5oJCWGRT+Z4o+gis5Z8rNw9qZkEUb1qmdJROb9O7qlRZNK9R
+NOo03kVvyVYwe/wgd34U2lbpBlmNeoW2dT4hUdod/rfPfnN/AZRNvrlcxYavj5tuym0POcgGOKD
TZe9JI4B0p8JUHDckyjLArGpT91pUS7ecYDRC9Pi1Erl38S1hyOaoBdm8SlTQj3sDujl5vHA63TY
YIczQyFv4n8Xby2oNhMPKednc3WtVsrOq02eXvutZs3K2h1IeCLqqk3I1CUXCMt/eLdheZ4XY2av
vHqUmOsWjGvIND0F7DuGnbjwO1JHrFKCLI6hUDxW2QeeKpptL0BPPbjZ4/3u5eyu9B/0Omvckvyi
gxVGqyFG94nNjO0pXBm8Z7euqA6lLWaTjvQZ5BfjEHvZ6WunCndcxauhUqZOkc4j21J4px0utg6Y
qHjmkrf8nM/PgbBQWPeO2H+sxlTn0lmzMS//Z1adjJqxz1IDmLHPnmSQ48PxrCG+oj9lmpRos3Ch
uiHu4a12vKlFy/vL9yPkaE2QgFwqho47miq9QCZX+WCVUu5mlsxrmYf/E2j1c1Rtr4iVJmPDBeZR
L8D5YHH0dQJ+vCgKbZNUwM0hZKNuGi2OsoI0JAD4Ka5sxYn3iC1di0aF5sdliuYlAvAF03l+F5Nt
oPnstffQnwY6cePcAldEyGDHyXdtQEuBT5VD/591jQijdtU0nrxrtqcAbutR3O59wdm89r+gJI1R
K7kJASuG8wH7i4gPjuhqiaeJkL870RnfNWtJogVb1p1ME/FHI6h7nKjdo/4TV0bWB55J+z68pqs7
oGeZBCWJ75U5kMmU3sPYqNlS9qVWazXHITzOYFh/jfkn9+yOeO7AamR04HHlNjQzVMemcVTgIR/j
G4ZTRfzZDQOiqZJHru/uPhfX7ij1gABez7AsloKfONE6CPh0sPp3pgm7kLSK1GMTwhgQfXVIik7i
o+VjnAzV+0sL19AXrosPumJ+ngs0kUW3tMdtn009tRSmYn50uLsVuoKdipOId36SdH4ncUiVWgGy
oRzxIC82wvSMBrwm/Rx4zm6alkGpdeQ0oWWTeo7pPOyrOmED4nqKLqROBrrq8GOSQmK97L/CNUrf
KOya34ez0luaBlyVP9onBWCu/6tVAXYPHXrdrFa3q3fCmvXMl3S+gBhbIqFokRGLalqcHAJ9N6dg
HUlWunyWehllzjg2GoLlamHRqqJMC3T0ugOv7IOSWhmC2X0x/f1D4ikluVM3RWqoNEpxOvvKmA5x
NRWgfsOtbdxug4Rwr1Cz2FwoyYWSMz59HdPXK8caF3wFBD0iSedRu8Yt9Q5Y+/DlMIauaV52XdNH
cOQziS39uA/XKZVJ81vTJJoWS2CMMqe8Af6vgDjDfYhR4z+B/USBwpypLNyakQaq3xcvWmtyrGWa
kiuJAT7K//sR5qFR/nt9344VIaSpSzVNkeV2uBiLvlsS3bCX8XEzu0NG+gpbMTRhUeRkUF0a/z4t
U0sVtvUOPZdnAGuwdpP+3JOxb7lD7sDiqT1OA1ZB0SkEzctjHCf/UYwhIVIU1C8GBgL9QfUyADyL
YJrQt3grD6tuTAehux6+tqItYjMVsmzoH5uE4nSWJuZX01uQKq8dcACau1sf3UP/eaUrFhxDuQld
9uuf+n/hf7nkoCjbGoIyNM40Cc90vlIMcvLuPJFZ/cPA0kyniUmI2Lda9hGLh015yhCO9aG2xV4b
godztmzjG6bTsPGBoS2JASvhhHzP904TYyMxSYfHRextHamxOy38BwOgsgKXqBBIMoX/QTqolmt7
CZMRhsj0gSEYlvCsoiPg+qZ5PKrsLTkWxLqmNnmd2gBcnEmda1P+SCQQu3wY36Hl4HgOOeVeupW6
4Z1RwTaHLZdVs1k2E/yeRql//ZcADHVEhRLL5wPD3GsgXi4cUEFtcPLaGD8CiE9xzDYKAF7sjZEQ
XyH/8Ologp4yxDPdt/CiyRjbYfWz4G5l7m9N4GTDjqbFmp9912pK884rxdIwigJWz38RV0fQqak9
3TUfvAOdR82V/dTi4bndlMPQbz3RTeI0jPH98I77dWKHXt+asKCY2vklmTUsmsnKqiVG3KV555fJ
cPG4ELWSXiV1ML6JEyOF3V8EzzmBx/0cO3xJMlbT0RQlxU4tQIZIREAIkEvGEDw4FbL6knemRN/9
wG9mWvLD5PFQPlt0lb5NSoLdoSe95qtxH30Zqt/VFkvex6et8Hn8SUdPosPju+WU2UEdOvTt779S
SkBfDCXiW3D/ve9bVsHgFWA71UANu7GF8idz+3rldXwR7wysTMQyEyxC4S5Q5+VojWR9m7NlEXxG
ZCHMzU0YKiLub5RH6jMPlB+W0CwK/jeh4j6XwD/C4SPoGhOxqSGoJ8Hu89SE+614CWBv73O+I220
6CxD9DhZe/rF/WpiDNWu4OC9lva/O9ZjH9Q0P85LfhXymh1pROwkrY5QRr4v3YOPE2+gWSsWrZ/G
hNTK5NAjcuZ2A9bSV3f3MPqfPW8A3pOWHff2f6fVhDuebn4wvTj5OeoN5p00LC5hhQs4GrJ/SasX
W8wzbohLGH0EjCRNUpDIBaRIFEXx+8ZXdYwbxD2fFgRrXNL1249MIyIDOcB6AjwPr+TGwj4GJnIx
MxHdvPDa49DQe6wmNZu2cfLs+K8X7UhzGBCrv+574IHkZZTe9EI5+zeeKanwB7IaIALE+NBMdQ0M
JumPpHWeLBQP0YCswUImcsLLlaSi5lQvQyB7rqv890t3RJrWFULmq9x1LbGJfd6bi6ETsZLhBYZr
gVHjwxUNALBU0B4x+Rnx1eR7+sKQm6NUMkMYRfNho3zyJiuRvv3Ep/nBX4SS9r+n3Qp8i7/I672o
oFByNmUWGVaXagQyX+oMPu1ovge75H9TAZFSRRqQPrwFeggzqiFDg+EODGDkSs1pU+1B1uqmwkSl
aLYnxayxDRNKfyllxnH4+x6uPiptqOQvpAZ++C4qbbTtKLtPk9JesQZs9IXigxv9Kj+cl2EtnzAB
HJ+bxNmYEjpJwNqtnJhGJhz7JgVlpd4YsiW7M1dceRSCVcMB7UaOSHrxvwLknCkkNNIg9EdG21c2
Kf9Ui8wEkMpQem1joZ36md1ce04KqGnhlC8u8a/y1Hy/NrmoSKZSywGiZMfQl2IToIb18jrXBqAF
cj2V63lfCvnrGPxyb6e+g62Yz4MLfTtu0H9hbLANenZg+GDf9J+WGcVIEGhYf1wTGXyyvEI0kkcV
XZboXIYXvOGHUqBvrbKiyTnYuz2cDX16Bw+ZR2D4U3HuDitUSP1C9nUGzvSIhH/NOxQYbSaiFCCN
6INNA3fzz4JxHe5touL6CDie8DVd5Y9pxKA4zK7vUEPD+x3VbAWIF8pYGpyohApPhlLlNkVLnWUU
h1fESyygu+PyDkgpJUvL5KZx84AGETsdHq9+2unL/ya9n3BeYW4pSZhp0az8Mbp8WyhZ0PsCQpkN
z3BA/Z8dDwSlbgonTilEz8bu4QoUglR08AuR2fkYUWLYD5DRhJhR+QWFRaWedgYevoyWNp6qvLth
Sxg05mbGY2xNTDrPcx1z27OIgOsHBU7+3IFfyE8eUzX38yQPyVI9oD1DiewKoYoKo3k6ZAtWHuFB
H5qYwlyonA+15ii1zOVYa61agXmsVrKQH8+vjH30TkoJPbvcU7p9k7n/nVNjYG8KFRK3XLsMl3l4
30KLSe3PeTG60S2pMMkj9o+rOYQ47VV/Jg1aBKLucVR+BC0l97Lbs+F7AMDSkcLnXy1WrutjDkAx
wuui1YMQy82FzfGxhuep0rlkQP5WsWSYLYDzw8ZZlhDKSrWYd2lr7vOWhgUjMv4nrx50vYdhmxD2
nHgJXZczoF3XRjAlt4yXpTOfVazxbBz0xcW7SlhEkym2YJXqt/ygS7Nuk6cYqy68XUB6TGfxNuro
C883zAlJ/i554sXJ61Ns1/TeqoTrqFQUdrFdndxBjMAVbdsjLa3pp6Cr3L6oo3L0TplpJ/a3Mi5b
gtoO3v/0LCDGVGQi0R/1LN0y2/aqk3Vrn5Q4wy9o7Cj8rhsI0gmfvdKm99yVoUi/zfd3Sb+rnmf6
OEcEkE0TcR/2/7DdrhTW4fHOYbsYg5BU5SzxR6NZ3uXndI4R+V28yIP1uz+N+/Oeexr8nFdvRALH
C+yTOG4t9O2ErCLOFWlmfEPvtmBrYDCSexPp4oFKoMZATLKcbd2hpXu8qqCca8DcFnTGW3+zEoMC
xG+92XTFnzwa1yva/1UVubPK7UZkopRs0JXVCVUDgMDLT3xlf7GPRBQ3e49n7tIK7lhm1z/Wfhcc
Jd4XwQmnUCZVzui3oYAPb3zetEkajJ6XdAEdua9kB06UjUVk6lw/FIUEv9u14iy6xoLZSOElJ7iP
Gc8PikgEPqRPWduPAV4QwqOleAQoXzQ8Lb59wxQkRLQUqFnOr9u0OWn5WiOsdfuC/jMU6nDfcF0r
B8AUQQka1fdFQut4X/qurlpmc3JwRLhCpJjmzKFVZv4mc9ilCi+FRE0CNk/J6mjGpZh/wt3C7One
RzwjDVa89D0r/V9gnuFtF7RDGinQ1eFMVCUxT4CUia/l6wkP9sOqhL6RzCPFyhH9iueNnAlPGDAv
HYgnVBe1K6VaT2dk75d6J1wkbCOnHiI2eibm+02ErnTA+1kxlOK8FQvXI4H9thrRmots51nvAODQ
HX1GgFqOki2WILdEozW7rYN4GjibY88Wrj+csxl842wEVG2O3rTUplsUCQ7XWqAnjMps9aj1sVSg
iBKcobXnyQF4o4TmrjYP8BKXbGYNW2gBQPxs02vP9LSEPXQyaJSTcO9TBT2gxCTA4SJUmu+StNCW
oOKxJTu6ksDkyWTVN9TDm9yDppb25tEdKWLvzwwTo4grIvQnFXFjx2dMDk0AgSYt5zTFoI1a4ZVg
L6pG75OrYXfMQtIovyFf0UEanONkGYoG5h9k+yZUk+SSHPbbtJNEDxXVaK4tdtIOK1nWvZu+1kTX
IRaBx1WEy0/vK8ucfBKO1KWeaqmLKpLlWRpHGwiIxEYk6IOC49UaLvbHK5vsvaux1gy4tJzHIhQ1
O/duJ62HsEFHZrgHYf+4ycvsV7lpRodqjubBTFKna+wxsFQUoCtkGhC4GqNiZ/mVWih1FVtovgRe
biKKU59gOiyJ2ntfk+Pr1L7Pf0XS2VcGgt8976Oqu3n/B0eYSwOIQLvQ88lXpmCi1asPF5PxqYqV
RDHCYNZy1XXH2aLnErwMzQutKqbnXHh/yz/9Adlp40mMkcO4jFf0QAH3CycdPyDa3C48/X0v0310
gZnHyxxHSOpMb1qRbBzEuqi7cPebwTHcdmvvNgtHWkM+XfzqbNvou7ql8WlyTUOJSDq0Rsa68OWg
MCLvvHgmk6OSoBWZUjPftOPz1OoOqaglsoCpk+12wkgMAShtfy4aLjTCSDB2G4bhxjFaEMAgGZUl
yyU8X4hhWuq1C0V4cVhBgUU0UXqAYlCsooPBoYFzx4cA+wi0G0c2ccS7ppOKCyetLz4Gcq97akOh
J3Xbehtj+1m4W24MZ88XVnJnTM1MS/LGFKwZ5bOZgERd/1x5Ws1eh00heJpeZa01wXuKLK/at6Ik
RhHqcLpH6RwQs0o4Y0OX/FtHeq5avPc94KJk80x7T6o0wltb/7LrmdsCvWDNqsWhuGWY1crzXsJy
weNCEgBt8wZhVQbY14B9ECbcGaiyyquO7ByPHC6FOT/CFl3jyaP5m4sbC3VkCDR/g/FDuZK7wBIu
lUJrxRD8znZQnKHbbRkJjRnfQI7HIwebrwccZsgpUeSU0MNVJpJVmDYfwlg0CkvClVIXGhVEpW3R
t+UcNjPDmsjTbW38CKGM6qFH/Wwsg4+c5cOVYQEWWRgMUMGRyBx+ezL1RCpcJLucVYmpMNjgBaM8
Y2c7G9DC5lkGfmBfptxw5Bn574GNkjJJvMVpcQv06c5XfzPcTFFGRpEQmA0zPo+BUfOo9E9/sXSo
pKthvliCGOJ8VwOObKkkUh3+r+QuLisIgFVdk4yAvzeyBn4viXgm7BgYexFXRcs9oDVtmDpkuRkS
zr9RgcNzX3bxxJEFUkdMgZgZmIhJ3oHLzPjJ1nHxs8/iJww2fcL4pHnu0VgI+Ky8MR8pH06tU6fm
ZqTCGIJee0p5Z1p9+IA+MD9pwlnxg71OyhKeocsE6Htrt7HjGLh6RD1mEpxn9bGhhVepLHfcwMgk
Q8TjRrQwJSbSBFo+P0nu0h8/A+Axuj56MQQc+ov7nHZuOvUk1uBjnECW2hQWLf7bNBNpi98vuTge
pAS5vNFHsJ6h721+YZrcb4rFX5wn45HqT9iwJFKK2mVZuzbc2a6QSxkXazHaHNvZUgtV9cqNLYOx
hr/Sn2p3gydnFQEQrggo0fFMvl6Nv8AvInj0ARLhMGlTx5KZqQMomjXK6RQLFJTgG0NDtf+04ywX
kSXiCdSRiC0KtV+SfvXB1pb4Z3na9yeklJ2po/K5YJV3nG4LdJY3NnvWQF/6iC4PKRJSF3jjwc8Z
x2wm6z2MkmqTJpquOiSKGyTxl9zRUWymWW7uUb3xhLoSawd26QjzYfltKFsODoTDBejfbnxyuOsi
R+M3qQxW3/seh7ANJLHOFS8LG9z7tQGkmbgQwIE4AAj6L2/m4sarMG8PzmN6tAZXj8UxzaG0R/j1
dBNzQ111ki0UBCBaewpEpjam3XL5wq81/uKptV5xuorTQeDZeEVWEWa2N5YzatbVXFIac9CkuUnV
0xhRwQYii6PRSmTQcPp1JwnnI82wBRH3T7vlMOIvt5GO1Om6I0bNQaN/gqt74UBshBj2HHLfwQ5x
NqXuXzZ0f90yExC/1qkIGv09dXMGUIMT08m0iVo2cpWKOkUQVH/RoqHi2+Jw9HQrB0jH+Au5SjYH
27Ondjq8tdxZLxe91q1N2/B+2RZsb2wdWUamPQZU3CS0Vye2sDbw/0TLc4mvrYQP9sQUUGNZ6R7G
Ozlorz4BNYijnvKAOULYLSliN6hqmFG8Q2oxJY5r1vE3Tyt+POGBPagE5Duf/Zl13WRcpgl7aMEp
xHe5ruo4v8xPD5o0svLsKJmNl6Ryc71ItJpWAAf4Q9zRibmPeDoFXcU8CKzdWsNFmM/OCQ7sprO3
vI0be2+3QxQjHYjPcFz9AKUpxtv8VYKKDIUI8+WjkvmuPWacGE4qmT734tppPraVZVuK0aHJeejj
vHbaX+amY20S8BxTtZMg0NY8dRHio/X7uhDGrY16jknkfMOBnIT5E2yyuafyq7Ez+s2flxZu6z4F
Akd8R9OMWXMArJSVZGLBstn461iVFpMY6GvoEe/XAARtxOtqyN1w0syJ1nIZLJYL9BUN2YU76qQ0
HPfMaU7UwKvN0i9KvZvCigmiN/2jJ3Mju+l2v5iqJhnoZgazN7JP9TS31OIpcBMaxSC5tzuazWeQ
d0JWElWJNNkZH1iEF8IVmsetuZX0df9bwIUbQMddE1gFvkzT2nMVF3N6Mvn7Eb8Yx2ol8zAZfTcW
w6tERep28Ws4bdcFxnoGRWBSFsh3++0p4ZtBA5IBdOs+eXsG0Dg0yo3fKqyFTJtqkc0gLSjTfa4o
7uPmMX+oBk2Ckip2Z2z5/UEtzAR1e5/oQgWbm6fgvvk4SP8SrDK1IDUt1q/1DQz4V1qkiqZNIzn3
I5P5Lj+6RTdwSa7NBFtKbD+f/i13uqC25RgKYYY2Jj5roUEwXa5OS9B5kNyl6xKt0waDt8nckj+7
h5v77nAwGu/WOk5LGlf71x5UuXYSARWl59reCcG7ZD0qb2t4FhujMMBzih3MNvXTKwERNcWuKvqK
Kqk8+P5P+wKDFuPLCNT3vCQfbPPwTBE1o0698TtQu+0guFkrnZdmQOP7dd40oKkrhYQeLjBiwOVD
f9NK8djBgbRchLyCFoTZgHWxLADKMW4/Q8yCxt+zkAWP6+KQSxLPPGhb9DHGlnRGeyj+H5E0ku20
zurLtpsMck8M64Wp6RCEKWMqbqO4AzYjY6MvMtzrGoMzWN8lCOwPnVR9o0yAPtyBfeTgJyrrIyUP
QfGusxk4ReEqA9jsvnRcQLZIHqedD2y0QlwzmyI+KYCCEi7/CyDlnlFsgpOOUplwlg2KlXf6oG92
3Qbi9LP+Pn+B/APt2wHIHrahxK5o/zkxcNaLkeHccqJ8MB1nVcyiwPk1Zulu9IVCtfW3vrvF+lhN
j7YyW6klnl5GQLpEE9UIAI2weqnE1aBTWYQpyZUHD+rVZZuKGSwFg9rI3UlYlj1zipvHP5hD78u0
5WvbgHYl23Oi4k4Re0i0PTNQ2Px5fYdko/mYcCMpecKXtXF9fgM+Kkc2A8ZzENdMCNoEPwnz3kKo
iL6pnnCwQ0H9pGT1A0sljULmvS3QDPAgJrSnBDm9TI6PjVOPm7e4YtF5SXJZtDmroxDlShwNv7n/
+67LSpMwSflkXAaPP+Sivk0nZSVvlxtTY6SQgHmX/B41YAzp3XmslPU0545/xVtyYKcscdV8Xqah
MHPnfcWytnzBknoIMkLMjZN/+frXcAnTeJWfv0OoO1PaAfHPQYoEvDbYwk6QKzRKWC/T1K1PNpjj
upsCMw3OV4x7Gui5HXQje5Dlj+ypGSbU7ihjEL7YYGfrUuykYu4mgeskMlVcwO2djrwFnqq5FeWv
j6dhaqenNezc+a+TUkK5ZFe179eI/KWR0+We2DU0pQpIQLf/+oyWKT/qcDNE8RyyM0iFGND0In9U
u1uunYN3mvpeusXDZSZCqOFmRMpHb42dJpIhNOwnqZNobkXsoIMP1Q7VdxNsmOswuI+SmcW/efgo
P7tOqzOTItWYsgtJYqKMV+86XU4VxdFMaouo3rqTgUk2sV+lq88qyEgFmoDxMw0UmwMCV6HY3v+w
bpPs4/bDQ1q9UBmKFHNDn8IF8RlJ/xYW9FcxMrvEhVxgfvXFy03628MILH7808UzU3Z/dZA/nxYZ
R4rDEcTkeT4QI34RaGV84ewWtEAjuZ1g+SvOv0Iiq415xDhIZSlSSXBb8EMyGeV7tDrnmbeez9JC
Ooqt+c3KdupQlaJEIOW4TknQnk7gm5NMPCOmJ8Cw8rAQ9a2X5CVSuTFxVZVyYUOR0i4j0m4/ruiH
EQ/pev4SajWLOxnfv/Q2W6PmWT4y6+osCU0ZyrtNZnyhPKu1KpYrTfNi4I8qj6cHWxVCOHGqTKqT
/9IqWjrAcyTxDIH5/uQ2NINyvdd5MgQj5eriI8g3HBT5ll4e0laoICh/Gw6GQqps2lnMbehYxyfQ
w+L4UkWfy26ppWz6kGMyBqTEwKxr3Urc+/wYhai/LE+DPVK8/WE4Ae9K+xgHQsda+VEw8gVr95UG
Vbes/LXMxUSZ43XvSNGyrgvJqYLdCIQQD3iRSjWfL1aYrfujF0ZUOJe22TjeCrbO10uqfLWVD266
CxZvrdAfWu/m63udoI3vj95LE/L34Lr6eCaDs605bsJpM+gtKlsk9e0HsAFjwsFjNW9XHSTUvqLl
vk3lA0EOlxrMP2cX/Yjwqw5f0mmDKjWjVNCXlXpi184cRVEc8gGPSJlGS1EM+Le8dZ2ShgweDrK0
cx1Kv/bFOzLkRxyeWLRY21FhcoLB7J264JfUZPVNpAHrcLWPAshVNHYBygiVH/gewKqm8Pp6ixWi
uQ52C7UX2T1wNSbUztl5phZDMvChiJv6s+j17HXn8JPU4eySm0fhwJnAp/qgUzcWgjjXFNySTBE9
TwFFgUnsLeb16/jcO2deiAywwE4mp7U4M64+blJ5JQorOdQ4vOsnlbhP65TX7v85UBrlOClGpH/m
XAD76qhCKO0Cl1vss50IQhJAhhU82AkQ+GooJ5A0hqxP633sYuxWUTYQ1LFWAAo+Qbwrll8fuhAF
/x9vl3bEFRelqpr3r/7aiPfAf3H7gtcFq/0nj8i9J+PgNeZN7tar0us8tyhIcSjPZHw266rYRpr4
OKpLl6EpS4W8Vi5PI6Wil4NPt9yz3p4aI4WhY+s2c5NZSkov7lHcnIhkUCo7rAfV/534K3Ysh1ID
TW/RxLAswpsLDMFHkmSJzkTVkqlasT87ykLWta88mGH1fWcRZKIliHI8yeM4M+5B5RIRr6Rmt+RX
UbC0tHoiwKJ+8R34LEYTE8pjg7oh01oYZQV2sUrkgMILTukdjfmUMwetpbIl/GDl3P440xTDlriu
j2oIQ1684/RHr6M/WoGIGHnadr8PLitOFIRatYYL4WN82h5REXnqAQBfiWbNkwdykl+rBxBhLpW+
/lFJmOEnkVn6IQsXK19ocjiGaMEMxNBLtMD6xIuM25zCl3p/orW++UpuVr6lPEiiI1CF4l9GS6Mq
VRD6WCgL8AYM05zVKuDDF1aa0lXz6PdFMEPAIfTeFFJK9yIzUm1Y0Q1CD5kDCGn3xr5MmHvd1xp5
e8FSMGcwOwBiTZHFJI4Eq1mJyoMDArJLpU89jLfcjepj03Otf4Q1B5p4GInMvbqrM9OwpuAPtm8S
3aF3e+7Vcb7lZ8Pnd4oiKWcX2I1Kon5+O/FWaq018G2kTqiC19ZIJpbd9Jjz9N9lr7knWkroE1ee
YMUvrrTvuOwChlXVGHjbL34tgDYbguojwEqr8K4EEXP9KmzrxXrwcJgTv70V8NBEodGJu4CZel8r
6jWsRPvKNFk0EbsStxOnwrZFEAFgIRFqfxZLBYX9rnte06yjghOUKZDLPUex0gwezzfO6kX2NLL4
OFd8gWoRm93qyeF24AQ/fputhHNq+rfyLtSqzFE3tF/SbMz1vxknI0XK5HvrlFn0KiCZc0XZJ9o1
8w2HpaHnjpXXgMlWNMMZFCPRzEqO8rwi3Z6OmblJGn9UEP991iwGL2/KCPr1bJyZ7WOuUGUKeFk0
sb8dl+0aksUUK98BtOnpKn9MSjGggx2iqjAqGionimj+DAi8OtUqzR0lxn5VrumOyAobocsga71S
M83SkJu8eFUWi3e40zjIl14LYkGrLpIwRJQS89SkkkP+0CMLLbH0vO8YEIdUIfg41hOJq30OMLt7
yKVGOttSydnfVV4VYxupy7J4Ie8WBEqOSDrtDGPR/m2WZt9gzHhb5Ze3EUgnoa4C22zqs5i1O6B3
dA+Woj1S2WJ2j++2DSdF+RDZMpfJs8jfuNUoYBVikm0UZA/b0WJbV5R4GKBsyaT7+E9gtrFDxr9y
DSZ+d58HHoYRfZ+rovEedFUA2MYKCWTdaa2Por/hBfROTE0GnldRYqJDmUoBFyVaTSLFLA2ZiZgv
P9dXdPEL8zxvz+f+TkBkWNF8sDalcrAv07L+Zw/TJ2m/2TR3AuB3+hWPVZzXjsFcFIkj4pS4lvaF
E1R+61etjgAy6jdi7mddk/mbAGuaq6wlCj426hVDTM9w460UJcg4EWW5yOLWecghe97ecFKK3wj3
diKKQi46d3mxuRigqI3a8/ja2Uff0c+fSyRmzukKzIXlCSvTL7m+Vm+T88LH96qiDfBWqs1NmA5X
K9SLRqmysxUvqH2mo4dkecbRnd7qE5sBYWoeLwtwtlQo7ZGQ5d9rdEIk0W2nbBPugAruvOgb4yDz
dOT57J4P+lPrq5xT93DhjEzZED1xAFzhrC0CXhnA3AP48eWb8bLHyGjamYo4H3qzaPecy3pSOSIQ
wbrMwwCjMdhyEmP64QmcOk80LwvRY2fwO8I0nv2mfjwZ2W8nR7pwAMYMMZj9L7YrDFYdxVstgbII
mSxfLYWBuyQZQNr0NkuIVWq3J+z4nndz/JYLMj0elD02lD3bU6zIXh5pQ23ETGBElLVkk8gTsAmY
J3qbqsX4Wx0KFO9G1yITWg7ooBLm0rm0RE1MB0Rcio0sNIOHHicCJpvIEM8o3RJpelC5dBcDS1gB
sItspiI0XYJTzGn63LbGLp1WMIZmdCUbJyPHC31LrZYqJKj1G63zOLUDnYH5E+fZw/pTsGi9fuYi
j+VMjuLIO18yiz3nvlvi+Ydr2RUxhMsaaWqxezLdyg0p6u4B3EW+nC9182ucNRnvOTWaVPJvVOPD
p5V2PjDfH1iBOz/igS72KH4wsOarpXCmvqf9C6C/2+QRkuZbvaIy5G8xordj4pKdYodb6mey4GGG
KmhwHxYcFXmVxswGHez9ekkspENuerWOZNrJiKiTrV/w6mup0guEpt6P+5ISMAkNoZRIs3tZ5C5u
Ov8pgZp7oZI45qrNDPKzLY+GAOqAPerwaSY2DPH7U8G1pen9MjQyiXJGSmoAzQfzzDs6JaU2P224
FD6H5419ov0L2cilkiE7E2l4X1rpKMCQmBzlHgj7Lmc+aMFVdVpbCHQ07jdcT8FW0zFZQfngUrQ8
O9/MdPGhFvKulC42lI5k11P8+NLyftC5rVfsx8Y+1mnPXRJ5/q5sXndHcFCZJsTTbOFGzGpQfFen
FO2Z+DklOu4AEeWXboNro7kSRQmIrmr38enIFpajjPXMRew35JxiG4k4Z/W/GWGNvEQ+TqAwFBTe
+0Jm7iKLxjScMmMN/WvtlrRWgONzr3YHCkdnNkDddMpA9IImqthjNeMdEI7mE0BGOUfECoBlQ1FL
yjawYQ6J7c/LuICdTCQvPB0t6jZPFyk5k1qzR2jP1+SzAN7ylZtIq9TK+x6Io254XpI7tCrTG+Hn
D+3Qw4UZAx29D0roDPsJU5pj/nBY322/eYSh3crA+Ak6PEtWstbv+zJqa4GJ6IQPeB1AxF+2/+2a
YgAjhICOO2TrXLUuRAM+VKDPA6Li9Hrm63cxH6/JG6VvvuszV2SnZFZtIa+WZK2lKGIRv04YW6XP
C0TFIYEWb6sxUnrjiLrl5CkBVj52ABQ3PY89bdazwzKOTO1PLvy7jEA/BNWfrvJoTmBDbUvmnw3x
ZjST86yYInhlW/fX5dOMoyCcfahLZI0tH7jmN4HPklSobm7XsALo8unc3jdOEP4TJq1CdZGrEj/C
hZ9N8rNxP1dvXvbIOstJD7xZayTjmNYEZB7XERRWkG7/UzMvsnu3RkKgSW7QlYMj5ad2lYMapy3p
rPtVeuAao78frsjn3si1XSxh5e1WT8I0CR2OUYrBTUmN7OgkPRlu/0O7pwAHMqsJDrDgmF0IGGtt
gF/PkmJReecQKei3tSicuC9K0MhMkl8f+Nu0Zc/lBrGxCf+QZ7mcAxQh0u+OWcIzLzAPq/9ZEape
fbmqZHHcdznddLk2oqubrZbvcfGvdzeWRQZXNqjnZtDE1YcEJw3n1tOV5kQ7BFDZ9ANatYv3B6ze
wH6ebEu1zuGBrqOv8vtzwgL9IfbFWliWgnALihsjHFlOWaJ6pYlRN9RJTpOwTBmNQ9YCeS2AN2rN
Ppu+88hiIPzESosxPz0QI7s083XRWq7G2URztBJ1Ip1HyuTFEHWl6c/se56Hdn41oOOaGx838nTF
+MDLnvrjRazjzGtqJKbxC3IOKgT4VqqJEPELUah9ZOCK5b/T5yBxloZ3mHR0A5YWqju3ivRAsV0m
PkwI5RyPEzypjfVJDsdCwtBBtSHTg0a+gonmbwe6716OR5XZosjMG46C6VaMLJdkW+aFzOboSiIC
4IEKBJOC6YtTOMkzmIUPC2+A2hssVOyCfp7m9ly6KEOXv5vsyfDEfh+stkooQXULLL8kl9HO0n1o
0QKjmEEMdskmhgWUU+WEB3Gg28a/6m8jziVUfkt8K2wdgr95jPkJcobrWYXU/q2mbnU1c14EYTpb
aE03934T4A8NTm204Ywzs+Fgx5yokuVU1gHV17IArE0hOjsfNlYxFoS3xJf4izQHQpt5irmiMpKz
kGWhAj6OPvHgQ0urk8HRY4ytpJHgVv7ZUPNnnEmO8Cp0QHcEcj9tTJaFytwfG7oNx4YAYnG2w9ym
jnC3BiJUYuNZxwkbR3sbL3IuSG32zkQvJW8J1EU59jPTcTrMw05I+vsTmtPi2CfqgYzzAqn9K+04
q7tN7TUdu5smGLVtQpjbet9BG/IEA96qcVdHhTr8+LWdITBBKm4jQGTxkhy35y5f/fOWwADksL6D
AlY7h6CRFKZJ+/NcaiYv6skvh0G7MQn5H298F59LUSaABOC3RR1EhNuzqfbnqn+mSnuwhzzmWt6k
icAqPOjZlqqFHJyiwLrDteiP2jVIGAQTeqkVjxpbh5QbWqEz4VOkuZ+ABITgkst6WN7fC4tgRLo1
4pH3qztZJiXWBY2m+n9frEN/fvfRr+ZCVkCGp4eUBJNYI3CUlAjU50mW34OHY7hyk1SM7bigz3Ci
aR6/U2o3BpeYYqYH9pazPq0lbO/3ohkr9EAdHT5uL+snMxVtZiQU9FcRwEw2ktEpoK9YQRajooDc
GNhKc2hEvBPfN7ZdRwykjsURaYC2iGAyaNACzNEghyqRWEC5Y6Zx/YhhQ+/DOwGChTAayp6Q4GmP
bmY+bYaHBLfcqXTgFq1MzYsawx20ohc1qaUvSyLnXJ7ppjK8t0fiQZX78dj37QMeSABkscsldykh
bCyjbjDGuJxO98tSkP8CthLNORJTbgJU6gXPP/g9gIg6Zyap6R5JNWXH4XI2X2OadAR47IGtNA6w
H3KjKDbD4ylG9w4A9IW3qQtg/w07crvTUJxxFVVF7joV0zraJ98UQrrxj7CczDTPu8nN1GrSn6YW
l7+nitpDFDa4VNO+iyw//YHdCep31U6EYA38doDeE2b2lpnggXRC0N2GsXD2Uch3Mh4t9Q47oAjA
PlyofHYG9ohLm8wGo+OlOfdtVPQxwRH6WeRrPC/CxYW2gT12U/2wY4DV1SpFS9Syo0XkH8UW6zLd
wXId2kQbQX6X9yq3iiX0+dhBlHZRvthe4ZJLH07g0BozPJKFOLpOoK21gSRHVK5ddU4liIT0sU97
MFTBIOPvrNnV5AvLn8XqEzxqVh3/RPu25z5r+Ryn1WC1psCOZdkm5nhnpVIOdpXwYDk1yyKV6uqv
OIyj8AinUloi3VyZeIQOIgI5yQ3iz/zjbW98Hq3dMhjiC0H6GoG0k1TecUXpH9F+rXVN6jCfE0OL
dp65cc7NCn9Q0trlZrEVl90lNbN5eMmCxub4fn0GXTv5MlqrPwXXiJrjB+OyzmZlA3g9qZ+NiTfs
qiyS0Xl1/L1YWACEOURqaVI9j0Pgv1duJYUasq3+6BMvfU/KJAOEr8sMzaOLWBeZXck9BKbZT6LF
tbxdj9Z0hwjwMUwSLSaDFBi476vId3m874Xb+wV2r5yXo5u4xNIQm6EApc7k1/MPcVnCrArJNWoV
/TzrSg5nBt8MbdzU2Nz4McU6YO6k2xo4ggWEvj73GsCkwCzh3/ukl4vkLcb25gkr/OUaygiKsr/A
fvZT1MLWHQpu7ryJQOIb5vIc8ZrQ09uHY0JJ8aCd45O2dJjN1DtGxaZuByieyKeKzHbkrM9bgoTh
CJqKbnosi69wgsME3lgomezsOiYhbBoP9sxld0qaDOqSiTd/pyDnG/Ox0seR0NrsAupzcIJd29r2
hzKZPrMKE8WISNAZgUlARs+tjyfXuXrcfhrXzZLl/kVEDQ3laByQ9xPDKfPQDh9QCE5VAwIc4BJl
1OkKR7bYn918BUO15Y8s82cz4G42gHJk2f0K4tvGkrRiBL7r6858Xr+mFdGFhaSX+UOdoDHyngn2
dFEsBnPZtufD344NUcxxitBaBEk/B97adnBK//xGZ0VphW3tdEZaImJlBcNv1AElgpYbvAfVu9IF
9E/32BJqmfQAvwjT1GMGHW93gvO2ADj3XLfJGvQZJNFipwBysoQpYRerSUpLxNH8neP88RU1h0Ax
1RMiBEAGIJ/TICgIJLCH/k7pLVRMsDI9RrQiVxq2WWbb7dPcmrOxCstyAAH2JT5Vj/Y4EV0Xk9WI
kXHKmrG1wOkSucdBpNrNljfLXNVeGbYL/vY19E/SYYshxvhUBX4adkoVf+/D7+jHeUSnc6gGJYku
C8sTAspxkMCBcBm1Kqy+JE+7lNoDYNc+cVsaqLRf63kyxYmfLUKe2ZXljk62EUGddwCgtFVJtBvp
sU15oVG1LsEDOyl+VLR++xxT6Y4fTZ/tRhdaM0iClk0kV63YxRTXdVajek63x/oshmyirr5PMsRs
l0GW+yK3ih2Umd64nmlJP+98RC/FFKHD5IfPsfT83VRm6eoxWUkxjkrhk47NgQDeXsNdwXDbdelA
tnDpeZNzlnBIudZueUeeLAWTSX6/1wob91bJPlp4CVLP/9eTOfHDgqTGdkxpoXajawOqFJk02mLD
i1awyc3BsIGSwfhViYBdrf2Ap/PLYDcPRUPmaApLuUTlCtCyUT3MVoC/igrch7Lm1qzCsL11DzcB
3Q9D1jD/IVAc4RDWegvsrDI09ni3T5TEOhSufolxkKts8VI4Y4ToHJrfvDci+ROy1+7FUld15z0B
89gV4egjzxINul50xW7aXzzq+VcEH3QunRa1Uz/RLNmGqRx2I55PjS+bNafsyixkXtUFC5aeVDXC
HGGPz2T4hi1YcgPNr9DIC2J4OciczPddYxdTmyn/huE2+AWojoYmYoLDUBnvBinfpTGX9NUo+Xzw
4t970vdWMMv9T0LbLyWP4Swk3fhurf0H6TPUgFNQJ9Iw4hvyOrpUDwO7rLDxcj9dDrJ3/PpayekQ
jxBLGI72KUW4EDGfVgNuZ6nuQDTApELnvDQqfeWEMkLAdZ6BYiNhUrh4cQ4vO0fxowFT8eubDwQK
RO7WCYdCf8RsJOON3Mcfh4nl/Tn/ePfXuffM6WW/HejmW+o8rx94Hw2GjmX0ytNRDZZcYMyyESHv
F6J09HtqtuiWr4eaiTTOkajWB9gFwCL6+X4jHTCZIV2MUV6EHUlDx6TBUNPCjmF8fIO2KBZbt2e+
4eVUv6P2yvqjr0sr3Ya05hVtpwwBrd6abk9izEYrtiDP2h75yOJyRWEUkpqVQCpHY5VaQLxOXD4E
+J5xN6WqzqIb6yqDwOtHvMgYqcdxi7sQ1yRUASQ2EpkEsBgLbkb7emGlTlPrk1+f/TEVNVtLRhhL
yS8H/0kVTpa274llktZiYTwrS2pcILWML1E6n1tIgovsuy2iBNUZ6/54hYTUaipW0fxs3RjzMJwS
aepVJc8Qs9Sgoj7fIGdoGedHrxp4Awi52l31pFwq8CM/rb89ltovUoYCm+wlZbMtLhnaXIQOYi2r
S75O0lP5pRvD9osX4Lb6ZRQKDHR4M8TnCiNoA306aZeTfIy/XkgO54vld2otdq8eERVVk5SOGFK+
JcxkTee58hH0tSc4WA2iMnVai6Y8UAqzTRUif+L/KWdIUKdJWg+MWLXe1tn2TAxTkqFdP7UYlsHY
Kvzr/vLW+n7AMsr5mnOPyr/+cMUBEjagnjOYsuU4DVWwOfcfOf38yGmmhIz/L8qfRmWyqn7QuQV5
6lDOtNeFdpjv80CDX/zE3F4+gm5MlmVX8orzvUdZhB2CAIEFQPwkEwNlEK3Q7MU5bdmZGuc6qVF0
rfI2+UQyU/YbtLYzrz0uMGL+KRADax1480dFFyloq7Yqvw8NRrjVQ0o4AO3lT9ZrbgFr9ZTawvoa
6vUBcw+5KHyFVTqh1uSf3ZW8WSOtExJHqzL/gZEpWUTakzVd262jbedA2FWIbJkNnJ138x1hOTvJ
2p8Xc1dCTgFoG+MV/nY5MLQQqcYI/x8srVJkSo8udu+HcsUaUfnK7JdREYPPQ1FUzJAHbWc9CAgU
rrAWVtQ5L8FYYMT4nhdWQsBg14dI5U+EGpmJixA1I5MXH7Vogp1vGNUnXhJqwiHvxAkBkaeRXQku
BBRvZtzm6G3MeB+7uDeaSoanU0I0idbYjZw1cMo3ekDY/5AOpYKhxx2TWXxt0YGGy+2jYEKwMq54
URi96lhmQAuCwfRJc4tnrv79a8pb6dBRY0yxtwkFvCn0D2KwWAXbv5PmMqocn9ZxoR9MNB68smHz
mFg8sIquFjPQPXDstZYJoTPEOlKRdk0e/ZF2YdXBJjSvu8OgnJszX+4XKq0DfHVZp+ln5DyODOy2
TnwFW7Jb9rhZFZjNa5y53nZrFT1wsR9DT3t18SVeWcozJ77GGGb9IVBNBblA/QU82uaTyFEFTHZT
3jYDozJnLcxpoMGARZmhz5+WZrDewGOZgMxjtQ==
`pragma protect end_protected
