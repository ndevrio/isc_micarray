// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
RLVK8YXuD2eRTZ6bM4El1U63vf8orXxlKbc4dR7UOXAS0O5NAqZ3lHrgJ5Bu068t
MCuG94nEiHyT6zaoOUD4YtxHAUYj6J8uzxzzCADE1d+uwVC0gjcrfh2J6qazAsPV
aLZJ5tpBg+LkLIfqahWlqeOiii2zKdWaTjXaH7j5WbEJKOizkoQsEw==
//pragma protect end_key_block
//pragma protect digest_block
9CNyCXCDvTWD0ua86FQC5SChShg=
//pragma protect end_digest_block
//pragma protect data_block
fJuC8LXQUNcnsHdPlYKqUa0KmmhmhfRxoO5LQ8LSP/mSX6GMfzBY+INsUTWSxWgH
4m79wkTyza1TfBEe83wYqysmxlYP6GW4FZfRR0EWFdzbUXO2h93SIStwG2c8rgJT
uglLt3/Qxv7iu0yggBrLinjTY23G8yTBa3NjATJnysiT3PDMZPuYiHI5twNB/ieo
A3/cmDX+mAgpM8SlUA6m8NwJLXumup4kY90Ja2vT+bCd03JBWvv4IShGRf3inC3b
DDkSB7P7Dlk4sEPDfm+W9x+1VHJ2IsxAqx+f2MugZwusB8qcTZxZnPYbf0gfZXS1
eZny0Xp9DHUOPwztB4YPZhaPp7/9yk7b9QFFpVv/V4ati3/wEpzHgn7g5PIJjHQE
9kpuoBqYC+QIfVDzaB/J1E27MwMmq5fE2XRT8am1LiMTOqHaC2hmTWd04rtMpmSg
IeFLbjYBToNWiRE71OSGprBuPalxmfg2AIliIe2bSODWiWcOcPPNCLWCkvwJ8g8q
UqkI1nRfvHCe075kGtUenX+xnH1VBqw7qT7dnOK6vzcHj8rV3qqTI3Yx9/FxM5lD
BgUrtzx6UVQU0YuMYNT33WiwinWe1BdiACntWbMB/um/zDiXyJJcQvG0u0P9MAi2
mdbie3Uk+GX2V09vSbCeX3luFGNpfBcF8eklhvH6aZ2j4LubXZ6+QX8vcD+V5PCg
VwIs1SxGHIaZsRgQrnZbSVN0rveVItOHsV5t77Tcf14+xnhbSWQC1ghVaEYxYtiI
2GhzEtOmzC2B6kyFIKZV7IgYPCVFkDrrtLVwdn/TR+K+5OgTrz5iEtF0l2tBaHS/
6TgFAUMX8qdu+C6lm9qgDpiUBBAbvbXrYodnclSTS5Hg9gPk8VQHvNKQHF5GbQrz
erx9SiGBViun17+NIkZAy7g1FJw9N7o706hYwqS2wdL4DaqnnHCIB06f5qyc5bQ5
j1ynnUiirqCVg3CVapI7Ga71JCjRb3oaCQko8jPZ333ncBRzaAy/zKHBXT5OgCge
rjn0kP72WCi7owQw/k/N9+s5Wvzkl3K4xNRez0W2otsHWVw8mz4Vt0KaAl0rWJUc
F2vGPtrO2kv8f/px17/mCAhYmf0yYsWQ3DSQJU2tDwDrsbevy3YqdON641mDKrsW
alMqhVeYsfumbVeFPL+ONwyG4VAm11xpcDloz3+9HIHmBLS/dtpjj7DoZHf+UR7M
XJa7CyUOWHz+ubRTkQNak1S4ALpdEYb2K44vaSMFDUp3U+hPG+hmrnED7KFtsBG8
RRpRqFfBEk45rStt7W4z2bKFfMjdHU1e/JyIapqVFkCjpvtAHCElKMjCtjNyC7IM
7VCLXRMBKWZtU0/xm/g6mv4VNCKM4YyVenwHXpo38me9M0PwC6qon2ZzEDNN1QMQ
HWjmOQgf3mtqV04etEblg0rbmAGRshMdR8CVebaUN9sbdC71+hgWIQIhk2P05/+o
VQFCLIScf6TPnEnSghJWRB/gREDZVR40n/SgPuPVfAkw7rry2LcSVfYr09jm88lR
BBOdcZuH5UY7hsl5+MoxpDmIeG2iJvseDp0cIUhUwm39EDLVtQZ1DxuyZWpFt18b
PuLjEFcRjKdmRWytJBMTj89QmnINxpC0suhotjFQXi3SpJlBIIV0+3iMym/3oLIy
zyQoLkrOJ23qStppIawtFpcvOiv+PiVCkioCBeZw0BRJi6K1o5rWMBwZdjTjfYIZ
dQxWe5NyvSgSrh/WaRPjeBV5UF8dLfmOxD2imHOSEd8y2eYrVvsVTopdUF5RMsB+
Jl/cgPW3bp8g36ZbizK0fW5T3LvX6DRo0twXrVyC+WHJhEAkBzk/3IEyEU0kaJ2H
67K3RVSeGdJhzFFmWBQWBIPKySlVCigaqin/mnIm4BJrLqPALj80R3MT3oN8ptL4
q8jix8WLV6Zy49s/Xp1rzbaTH8PRM+0TBDmeW1YJXB8KHr8kZqpzEznuzFK6qLNQ
8dgKP21STXijdtoB/iig+hvAw4y88zgCM+9uGI3tL+dgxaEDsQQ0G3mKdegCFmDh
MId4meRxtAXbwK2j74n+QQTy+UiXoQIqE9LyJlsR1zs9qHELzeR9dLu3ZDWNNz63
8h49fhRegDYzF4BNjJ0amxpHA4qvtsnNWPCvrdGEMDeHY+hXt8cgXgG5V7vVEnQB
7sgRXqxj0Qbq4YZ4CdyimqbLnRG/ZXpd6lV7y0ZrBZ3ci+Z67kI+mZyW3lnESd2E
HaHvfxuyHqEkqtEtOu193SJmFKoO5aUDIMA1uZ84qCYDcujoKR/ZmRQ1ue+tODdX
ul+cPj8IrDi5va/THOw3BvNDMV9B7DwqsRPkaXkbhQLxNd6XzVyKhsk/BhkhoTyj
nSx3WJ+sgPu8NmQFileajC1JsDh472i2KWopwLKZN8HtlMVbBmQuJAOjdyOsOYGy
GtABX+z92VNrLBhJG2BD1TIuLkS3W4u2XgKGZM12z+XZldXm/k1iuD9rkTqCZaR7
adMSAo6F7LZIkrfqgokD6jOyJERL1azsteIbjOrIcoAZ8GwtZ8DM6QVQKIcN6glm
HgSKd/1hq2H9XYRvuwjFny1+73boHBlFDt5XN9JYa9guQmF52sQZiwFihRqnszra
BF6sQdCtnszgDLz0fckLRsvK7T5k7BfPf3VfoHxvV7b7t55cwEaKNYA5FxrUlVRS
JBN6t+h55RTrMWeylc1wt62q7+LJZWb4FZJ58HiJkGCkwpFgIlm2u/f9efMiYbVp
xgHkd9N89zEPZkRYq4dUhKSkXgGwJen8yv4Vf5rrg/cxFq4Ut2bI/NVtUbJasdua
UBI1NyTx1Qz0WiSBJzPOsHeI0caTle3fRj0eIm4g1VnqUYmYNuOUq5psi8rRDXWt
+H+QW0AjP/mFYog8ra4kL6+aoPDmOtMiWQ4AfAliymCGLlisgt4EE1fGbYlq2/ZK
AXSHBu93SrXNavavZFTu8CttolAuEgS/AhWPA9QZT4mhnh8Hzx/6lXEHm3YMO7/r
a59gVfU1pv5tl+ZGVZrm9R1TiouDRQzSO86g07qnCRDmI5al8KwuOJmZF6Ttn2rc
EFhQcg6hmtjrD4tp8zwidBdTJz9dog+ch7dgzKzT5hQzmJR3GPN5YIsmx9NCkX/P
qZ4Z816zhPfOq9eanWfj+Qaw1GiddWBZYqr8F/of805AHoqdjXQVnb24IGZCq0pE
N+oXjJWhII31nE917w6Lt4mgplLewPc4rNvJXPVn2UEsbQZ+8KMsIubXU4LcIClJ
/TPhG3zRbHwtAdARdax9/IbS0nVSJNdG1ulKvAIpLjKHHZ+koKAU04UTy8JN93pA
tV8l957TRuZGZCda72OLH7HqzDn07bZGNMPh1fjIWImUFVu1SVERUEX4jzdcWxXi
bEiQP7+1WbnsqUBQWD5UoNE9OOaVWsrq3seKm+XJUOwdsAY8bCa1C45Dk1P+lCbQ
gGYB5yhN6ICMUkPJrJeGt0Cj98EI28IFxWQl+gBU9V1YyfD3Byn4ZuPdJUaFh6EZ
AsORvjZeZPSg0Hc2D9G4NwVnJxIW+oFIUR929EdKE65jshn7nbQWPe8CBwfDT+Rd
tDIS/ZxNkQ8e7kavK9o0Rj3WxF363YeIEReaE68q6Khq49DWq2lGgmUxcgxpDhXa
MIZn8BrC9QnUKdkEFQqKvigp32iVATgWw58WFVhrwwkIq1wdBI8GulSCI1UNK+Y9
czsl8nhyEi8ggiK7iKr0UgpDR2tyF72VemmbpBpDXwVL1m/qBFvUby0K8tT1bdcd
ZhMbdRkpy5B0dglmZ8ywUGDHI1j80G7pFgdlV7XGlMkRTPv/X58zDyADzeK8h7GR
ifMONptOAJJzjXlry4UgQ4LDg1EK/6jVV8iOTjQH/UvqWiOwgrPRk8oHaBFE0AEH
Xw8bXbzAmMBISJrAC/pAcXypiuNR+axye3Hof3cwJJuYYzWTtLqQrw0NmPiUKvCL
fblB/d52w4XYhTIFXjYPkkPKzwRwv+FYSJ7aAl3/TRNleS7w+o/u2ep3z036fXBv
ivG0sdqSICEx7nsJat3ZwslMB3qzTugtf2PAgB/2lSGW4SlxSSzILyALj7TZH3cm
f9PKwoA5fDQy/8GVJ7WqfSOqq2/68w7p+zN72VStWYzYt/YRwX5jFF1EK0XL1HU0
GW5y7Cucn9nndF//BPGePYSE7S7T6/i/72ixms17c82AiRGjO3qrCkuVnkat3iN+
KDxDuaR7KAcCzSpFkYrfXqjjyL2lydfCGRb4R6D+0wEVTdFugJiQdQ6ejR4//qk5
rHWe8xddbnemfS0pxGw3oxFXUp7+jRp+dSy/IQsIF+VE5Q6pujzalJocwR1lP3s1
67M5zNQKMMCgSNATAoESIafqyxufMU3tIel7IvylVFd3Wuq7+ZW3fABJ/fRLITmR
ZdeyTeRQQ82uvQu9Fickvrb9dhfqohX3JGNxXOStI1xJxnYzEWcBEW3H0A++nIe3
SSmuAVNHcfidygxm1f/DRPu8JG2eon7qzecUPahLQqx4BbJBPwok8H0z8yD8QnRB
kAQY/80TtOMcx23g8nARZHJwkWtdJ0eSUTz2nOSo3Xfl6glSD1or9K1moayoEhlk
apvy8Njq+AGbh4y4NWVxYRXwr7ZyCEM+OE1qGdS9yWCg6DFPxkcp/q3J1o9nwRpd
2/OjFjG2lE97l9vQkHgv97Qglei0ZUQpaRJCizXnlXfaQVgmrzTc6GiTFai5Il+H
WCxx4fSaTW+4VX+2kwTWFxPEwgXz6VI0yEpPbQICYGPrs84aN4T+n0qmADXaNFbi
hhxACUTwbZLfPjC3bT/eYScdqNt83CjAMDgLq5LeiSVsoabwDlJGZmyE3xV2vNsM
i6KnCjOyskx9FuRnbp0kxPl1Bt/PbqUIp7TPQND6jDZvj9zP2oOCI7Q2ovVweB43
8Rx2RmLxYaZBIemhzpe+5Pjt7p9onNG+V7e/cqs8WmisvaIrFhUdpL5m+8eLsuP9
r80jDoVUg0pr59GtLVuYjtq/TJZF0vhdXF/l4JRPZLPppa6UBLnZLbXr1/jhiiZf
GogmSxwcXUqC0+lb7EOcmnwEFmfAKJrDe95qfOXtexYwl5ezC7xhXVXG5kUv/WVC
ybghKNSywcxn8WBNZIErnd/XNq00NxCPSAkGlVB5Fewke3haUSxoVjGfL1ePi4qI
7zORFa0ZWe3cIjHV/PKYMn083Ixo5yZicGkSxoojYNrHQ2GjgVt+VvHh3cUDyNew
v5CirpN+KzOIl6Yq7Gzc1sW4GMao0PqulALPCCCaf+owVMIguWZzzjHDfGW3Q+WJ
3nBTw8KG9PZw09/6wfPa3RtVm7dX2jJxdLlsymc+fQGyupupdD9+QrrUKMCxrcKD
EOD3lJ48BNC6eWT8pPLLdpQ/D+XfLD8jnelLi/2iNPA03EsH82PzI8fFJAz5Tlko
9Pwrg4OUZtvZ5v/84eLajUyJ4Ayt4WTL43Czn1wgHq9zj0E5yRQ2WijyDbInCl+I
FOCcsZ3G38gV5+9rLqq/leKDluf20rm1I5vaABLSpgM5opwljNf1JFvV33sVDBZ/
m8as5izwFjwB+yijgDeucIh8mf9zlf1l/mpmxce6hOQ1kh77mYhph1dDQgDZMWE4
P3vi/gE2Dm8Rgojqf9wDFfTfSqnc40l6EfO2DSf05HScl84RCGQwkDIvTZ0mo6EC
C4RQ0tu08xEXvdwYLJOn+lLMgL3QgMesFRBO07bLU95rqhYxzr6qAZ8F372LzQr+
m6MZcHh0GaH12CSXPOELN5h3WZCSxOEXgyl6iSSd34f1UUA9vIF+20ZDxIEbg6ti
ehLkBXHtS5OI8JKwp/h9Db27ZzFz2wqj2iHrnheP9AzWj4lUOMHPkUR7wYCg1iIg
6HzXgrH2yzX7XQYF5JuxPghX/KFvb363VwBHovz2PHmZ47Kw4cw/OCybfmx+Wn1C
XrWfTsvPPWczYZI/iPjYD7Q0ORZLysaOPaR6evl0NHbFWbmSklfTKQ771NDvqw7q
pScUwQ7S32zT7l7+xR5gwBGjLGwKSLr4w59ytdC98531Jhz8xfc6mOmgqQbkmHDh
x/50RODazDlpDI/d0M//Tf0xQrVU3DuISc+PNQO5X9Thf8GYYzp6sDhlzfSnsiXV
up6IaeGTRedY+BbVgvGjequrAeLJxVmG/1FWUOCH3l+rf+ZmksTxHBX8KJ08eBX5
WFiL/STCaSlycZgYaJ0b8ON+dg6gIdhzJIxa9hCFDm08H+DmQvbShvxryWowjzj8
tYBPtOBLjkjrrrk+P/BDEsbTiZL+kua1DHMU9xi/weRM6VRr6lL+vYMUpIrRD04a
Pag0zH6DJ7YkPdJdAcVBVAfNdq1aqS3KZ6pWeXCV+qDlZqjga//SHyOPtc6tMY89
d8sKK7IRA0mMPHEIJFghffv9Sdy0qDmvH7YIEgptp8LTnZ2uydagm42jR8Zwbiri
vTB8EmsR96ZIvZv9Fk96RqXm2p9l4KBIiSeNLbFxIht1beFCrtm6m7EZlEZAq2do
+B5thevnAWkt2rEvmNM0nesghzGAtJpBRVq9HhZWS6ugOFZuovam5h/F/oaqESWK
2ZGqN2VkaDLrH0Di+VJSYLf62r1wUY6+CvGw8CtsRfJ9APBrRSdsR6U91BEILo+2
T+sgbsDMRMfVMPmx6AKq+tiOvDyc2PCJP6UXxRU6/q1YDf+asaRmG9NVdzR3Fui/
rYgPUjac6qqkvI8cy50dUBChjtr6z7nvQ97WfLmr+HGMmw1z9Z4UF1bl1/93H1Jx
MLVbYlOWqVSgB5i5H4UZE0jk220ibTSwdo4NVOpfy/mIR7GjyY6Ay+2GG6aP8951
uw8F7yfFHGt7NockeOmzKbhwVjXv9eZ5G8qZLkhwfsmyV9UP1HIhSUhpw+/TafqB
ZCDChv8KlSHQfFoetNPkypQBZvWJCqakiBqEVFF6fnVKgWJ09Tjpe2Uptozjio7M
MNx+Adb+4o458YPxCDYjI3c0k7mMbOi//TOgv8UaqEu2VViJ/eGJLApwPm7RkTK7
vQeDFiYeJRqUxEIwgXvtuu6ff6NIoXv1vloggiqH66HCZGyi3Q3rbtzZgjP6RCpe
lf6wxKEJ+L8FQOhwoKf1uRgI0eQ+Gkz37aRHJutTi2qM5J3360IpyiJnIqH1P1nT
M7O7iJB7OCiVSY4xj9GuXMW4JOL7Fs3k2xriq9APNHtEKooNUkVUZ1DGctyu+Sng
mzVhjN2QUDusr3E2NFSY0q9mc/HGjf8vpu1ccVJ/PgWKQXgxxzNkwAoUgXBMLvJ/
Xowp/cSmuiAegBYYeYTpZu40XO+8FXhKOSlpxos/oL5U7tsyhHDn+R7y+lzU4t/8
6gOtQ53MnJRHThO0SbCECS3gbRekgoK9/BCGMqqAB57/LBXpJRkQA8hWXNbLDDBd
z9ZbcIJduvgRiPmPDYMUQArzK7X6ZtlUauT1hrFG1abG7+3fB9yEuUYljnly8mSk
3+G4glK0NygcSZjrXpdsMf+LUS+xu7Y9QqgPzZfmgxr9+Xao8/3CWJZRlvTlpDIr
4OHTXGaf9TV2dUs5F/0AmbeWoEyXKlDO6vdcnQFFyiDgRvyakXP45BLnyplTXa7Q
RPZaLtTPwhJP/0L7FatwJ6MJqrQLTJRE7ZgId6dY4p4w647BGqs02ltTLwpXc+5C
KOAsi25ESBpvvsaRI5B3NwSZldy1IUsWQmcb9/4fSacs2sxzUxZ/6wiRbkxCXtvb
GsaYThnGqBKGTSNH70OBrCOZFv0mxKmJE+uJ6x8imPTzG7i97u4dFvtkH3sCvm6v
9kj/6FE3KxiMyMwCV6Ai1l+7Y9WDNGMroL81FoWC4MapUdJhdOjGuK09xAo2FIhE
29xhsoqa3zHrzMxvnqOfnF7Y7dyKUyviyVWuVWLS13+FwZGRvk95wyk6b4dtLoBN
9clv3o58W/npaANBpK7rLvflnp8QsG74gxVgYYJcnnQCaGJimwOo1It/aQDLtYvk
/uh/Z4EuvKvKpArghHaeauOsL0CoZp6+DgEhkWS8fZuxPFcW6R1kpJ3E6m288cuP
xgGDnqsO1QUzKQQ+r2D8ixNbHrOhn/FbNoQ2twnc+g7IFBBMUkm4MXHA5kT5Kv0A
o2Ai9D5QaFrSCa4WywQE4eSXRW95Xd4st2Gc+DNt6+KzwjTAYDprvj7llJ0uCmZs
swOMSNXwxvtoZ++1UXttFXAz/1irFT3czwru4rJgp1edS/k1RCpk2Zhvfnvz2Xa0
1DLCg0lBrDmvFAn/VhdSueUS/Mf3ytMRPnLtlvAj7I5ltSysge/sdb35/kmDWuK6
WX7xP+qgQzRgW0buplI/K1R6vIfgFLBDYvZqrjRBV+vPysYIjtaq/5wqvoFSpYKK
8dOgfa97myfR8VLBOzwM+U95UMdXPD5AA57H1cMLmQX0gYGtg08K7wy9t5jo3h6S
gYrIeD6MnwqejpGIxYmht1XvfJsAylto+7h9Cm3xXQz2oilpZGf30sEXjQWUgQmg
rYQVosa24Qh9WmZ7cUcnpMIq9OgVVbE9rWIvNbw0u+3t/iPLtwSZJLKbf1gPh6QO
HylkH0IPMH8Qlfj5kFdcgqDcb3qCdkGXJ3rROlrGNtG78XX/Tvmp9TeGiebZTojp
g300zHBOwLewi++rbT+OGDDMANnQ8IyQo2YPTJrD0f9MZFJwoaMduXzgpiPLcAVz
Nbr0Q1TDy2n0Hck6T/d+PAfGufeU2/a12Rf3f9oEhxsdmoxYesStaPF27qki+Odw
8aQcA0BACO85zadWjuF53r8ZwNyRulKKX+yf9kuTk1x9OmyiijUK1X0TCGg3M+Z8
76wdZinr2e4Gz+Rrm1ekzGYrrBfL+49K7mat5bWne522zlOpmVQSZdml87NjLmOX
vr7PPIUXipx+ecLmL3Qzqc/uOr7N821HFrmYs49RHjtMQ3+f6eIDFNu4KFM1wArB
cHgpKFSg/bxk/cVP1oKWhiBq19+fP7wqPq1AKHb91ORjlvdfdY+inzFPn/9Y/7Z8
dOEqZT1+1LG5l+zwv5WM6BHA7JdiWGW1yvtwThVYFmkdLXS+wDHl1pKtei2pHdAj
SOQgA2I/8iG/r5Q9hdT5EpBg2YPT7rTD6lBFacN/jTNB2tzQflxhdQd4AAfJCQBY
VEtAWHI4ZKWp/mfalZpyu+RT+JcrI4Zd6xdUsZLkH10SLg+KHI2GBnRszxKjsJ+m
9vIYgzpByRELE7E2vMzbeQ/yUsMV6766ke5IQYGYvvvP2EaPQw71Mxg1aTQKpe1E
fw2XxOzE9Xfnnp+xN2ZJ09CmZwnKfVOoxPHxZ9X1m4QfXL94VDtoMbb22qz/7mTf
nwW8zY5mvub9S5oL9d7+lJvP/N/IC2OcsIZq5ep+iORWBEEtlQhDplDuDRpCdd5H
IxC2WFDTeFrIEE/qjAhNbYMtlKykkYDIPvAv7CklGNexrvPKxiY94hw5Cshr6Xvn
/TyQKfSkN84c+TA0xGgW6dIRjpsmmAYeQI9u7QBvnxm0L5yRL4alX5wIQaySTDzU
p2p4RLOCf54++/mNuS6pO8lzl8aGvm7zpw+tmQzyiAdd+xP+xjAjnvzFZGhW9wCf
TgKi+SfqLPyJwPGAe0i3ruLrdEgcyjDgD2gbWcVO4qBgg08ApC+wXsnaM0ha1xST
jAulFQZqQGXJoHJmBD3YYApgQSiEdMn5fp/4peLvGSFVxNoGik0Y9kdC+J5Sq70O
cMNWBWrK0Fc1xwDTWm0aW0xzyOnM8oSpoXCIWNAtZuPNRNIl84K6V0ByKle8gqi8
ppr27JNRE/81AIbo3qurov7yy7qMZJf9STmhTrMua8RG8YQ3SKZ1Sft3aZOR4Xx5
LzUbnjqeJsiL/SOvtL/lkLmCikx+CaTSOWz5oZEITR9eWT9wiFqaf64EgXGFxQGm
jk7E9OxhEkZGGuE0vT+mvAEL2hWzFzZYeESGmLKguv5I/SE7VNSpPMGtUmlVJaiw
DFYMCich1+cnWEWBvY7mAhrFqTAkB8m+FIBQOa+ebVTz12o/CexaqIapzJnPDSQ4
OftRE8+LhgCZgc5ASu3KCCEIrKBi+4Q6Tz9djkg6meBh9lFQktZaXovKT1YpNdHU
d6GSt08b0+2f183XkqryDJ0vjtA0WUI5653upjBZLB0itMV/eAc/KPe2fjIfkCW3
12AJOr0C0RU8xx9vgpndds3HE34hDNGubm3ZVPOIqma1VOYa5eJj53zb7ayH1J4B
Wam1I7829wu7aqVtd+/L40Jgd9/41epacljNpPtO2vWQ2TSjy9xZf5gaCJMwxxAB
dpQw59T2d66TownkyiiVUDNhe7j6N5eV7p02RKp8DQNcHvhx1LG1DRwQ2sWLyl+C
Zk+Pd393wAqJ8DEvyYOdJCxkn6rmHatigoAGsQVGQdUl6GDIAVHuQ+8RHFYUt+Op
DqAMnUu5pzruhesFc8fXryMYUd0UX6VJAegjHFIZNduY9vvvdsY9RVB7EUoa+pqB
a4mjio39G6pulgrT4eRT9JBhNkk1M4mcZPwkZM9vLZDQdZFzNy70tGLnmQhHO5FC
3SLINTr3QQfJtpkR/xQWT5BCB5P07qL4Y3EokFTNe/P8Vrgq3WybJovTB90OAUUg
huZgPmSFzRa+z5CgzRwi7vPj0EoUY1IpL4lnJ5p4pVQ5CQI8sFYI+OWhE1K50YDH
8TLvQKfjOltsfm/Tp3cmsvHjQFk45JpSJD9b472SeRF6YDV5Ye1QgPtHSOdWdv51
X/bwQXt2F3f+sklpVRlMQp+oe8zYT6Vb1FysnrRJuT7SXZ4MKKredeDRKW3vT6Zf
iGgJxgkD7d7ruYN+dL9yfIsFuFLDlfQiik8YKWm0ApFsqPXb/bmN/ukZAwaYcjY7
rm1GoOViGFvLxwB6jiKif/sgVTKN2HiwZpaePDirEC7tGSs2U/TX7A1hdptbCAXZ
AXrZL3bMQrSJVQA5jq+kuZUtO3490mlUt2WgWN+NF8r5zGadUECMjW0LXCBaTeYp
wMPf1s7uL8n/LT0tMXisOXW6IlnoZuV09pv7lSEJplcG2VOJ7xux1E1MS8AsB4pY
tFk0iAii2PhJPkXjwjqEAi5gogG2JRGIG0EeJLr2+0DFsPSDgs//Xg79P0O8yBMI
EgCi/K8l5CGS092wJFs0DKIMPywVd6LI2Y5uaHrha/zAp4c3OM5fn7CeMlcDFiRc
8yag7Jb+jEDX6kNcC6SkFFD5c39g8d0vxKV/hfhuK4ub10tkHJT4gVDmsby0aq8s
mQGkdjimC+MmZk8jnSWkv2Q+3GW8T7jcs+FeHz9mZAVCAvqA5TOGtm7MXMyeuVLf
c6xn0eZarInyCdAvsPmWPo3CisHax2mjOi9wDp9+SWkQupfx8afM0eLsxdwKfH1A
t4yOJNRhYmPBrgigprjlKDT/uVX7svLRQHMZKozAZPyDcaRpR4rHgAIfYjKVoTNY
LvqfGcR0ozuPiClVJeCdT+SXGQErcgegBaNjLYM+Cv/V3kiRlxdKaeHU4WJ+8R7q
qn64rFCj0qKC7its8h4QdWmpMbpht8QPTG7u/96e7AeinHplxVBoR0dgV7SWjKwi
KiNy+MNdg0LwRR++MfayopR9+TZE+ga0m5T126N9/Ls8HtpGqXObasvXUj+OYd5t
pJkAmeZrMZf/jOwD3WuHlRJNdeI4a5vp4LZtSRZmBjlBZyps3wMU8wCUljF4GLhr
0eWHcU7yKHZf6+ouTMfgFcZFarCKBgMo5eY21iChNTmYNJqpjb+XBgYSwXR/vgr5
QAyNaSNOGo5IkNmmXfGrAENdEQBswYwYV3Z30gSlpwbgXMDuBPB0MPTSgW5TxuDj
0kMNvCv/isWickPySXSWg9GZ94nY+ZWItK8/IHnFoUmkYmUnPciaPqMV5DmwJ5os
XC/A5B1NON0vIIWUTFcK04RUBNiwRO6hVSBneUh1pp6yz7uV2B/Xn4MQVB+yUpU4
D1eiTkJwXgQqTITTjRXwfmSEzQ0OUZ5YvNa9s/gR7FdorFpyVCiYX8yF27Q3HPPy
x3YxtWA6ng5N66y6B0D6SqR22mIiGOYqSA0gVOkdXdpAO+uRV+vk0L2+24XRWlQi
tFRcqUixo9SO1pdfwFm4mgnAXxVzZAGgxMhj4m8aFbKUyzmfyx9JJ1YPo9JE/IYI
xrTVBy6Ms8CCnOvK/G97PfLPfT5PMljSwfsTnF03Lq+Rq8UKVMRA7chLzyH3Y2KA
By6TNKYwchvWInuURl+Zp+59HSDpHcL9qb1uU/t/UetHhVe1F/3dEtDvZW5bceyK
UBONUYsMTouquFJDLC1hZ5VDNuwd6u4pTjqBXu6+UD4mk0G0eY7QDi0lxI2U/0Ea
pyVVLmzjQpfwlo4rZ0mlnSfWO850iCfJV5JtnpVAJCMLur86xfsSKgmR9amnWxGc
G8EkLMmjLbEcae5jtn/yihwWGuMQ9HHLzIRldYyL5Nqgy+o76jWssaQBRAzlsJkH
epcb3H4SmeRIZyhONhj7S/cSQ4XvIFZtDzfD43oSoyU1QUs24hTHY9mxUS11QI7G
IegyVCeGYg7KsI+LnGcpN8P2PFlWlrNC9IKh2341a/ChLvPgz9gkOoAYIuwpI+Hj
BHEA1EDJLwPV/VOKH5XczJzC21sfj7+KlWs44Yi9c0HZbAgbQT2ofbsBgwGnaRdB
vi+8fCrPaiwWnSpdFiQOodB0jIAmrl5ERnf/yeU8Hnagau9+G4Hjxzt3VzOmAtTB
Ta3Sqvck0eeQfHETV9z51BOY9zVPlV24OHo4KmC1zoEV4YeellClaqh2hfDpBnJn
ep1y1J1p3MVlu5T1QGvIchXbK7bfuOlUrBiTeJsI5w1CF6Kgwkhvjmj0znTJ0uj+
AMNFPRjqsMcmKrG14UyhR6SUpB4eHYIH7XRY41GLjSdq1ZBRqKELIS2/7i32ALXZ
hrryKsxl6pogrQ5Ue05Vg/5oDZTCQqYoplgMUDUnjZk2bS9UgTEUOYSTUGmJKahQ
s/wTBRqgx4TLeI69CJIXJArcVNwYcWe0u0yflbr2KO3bWKebqEHZTJ9nMFOU7rKD
SN97LRhk18FV6Zop7CYhtFaCDeLu1UN+NdzMDMm/+6Mf+0EPSJ9WsNW5J39Xq+W3
4RL+jawWZS+FiDBVwbLg7aeAnNyx4K/ckRN6FyJABuCIyNdoGEenmJmJwMf4YMO/
A458gm7dBcbXWw+AenOKJJXfmC1/rAAGNgw/K5wIOVdzRzs2umPLpWGudITleKE6
H96nPVBTjE/0/hGD6z8etl/BwaTZBnJMVKVAE1N/BGLCsvETjT2cmOaKYD4HqloB
cFWED+cz0TVyOxi7kXsdU3VIZh9evc3xPUpvXwc0Katmj9av7jjgbwzNcfuB9oZi
5rscJT1Jd+J9g6B5PG/NG8gPYp84H2lWpISxubFsvphb7TuMkUsregoUcL4QB7/8
qoaMa1cedEKrYNz9b4XRgUf6zcVtPWxQ1jLto9zWW3QGKUzQzZYON9J+NzauAlG5
t9MleWmbtNNM3iDL9yn8DLnFLumqczbbqjjThXM+yeHSQITT8jO7WkCyq/so9Ka8
q6zveObx3AiXCh3BDY57ay5cHNa1TRJBEypThr+s2GFxciRaVl55966fnaVtn8WF
EdMESnJ8pbNQUS1P9+38alLK0HAkWxRVJxlJUKaUWTYqpVqZSKqqKt5hZLV0BYoS
5CBJDM/qx0NrZSrJfVkpBPr4tqZvTLnRKHIkuS6sP8qQUOe57Wy+rcQPdFwyWosW
PMJ6pUDIMxtFaD8E4qWaLT/w8UZCoCVDwy0Q/4plIQRcGCyRO7InfA0sI0DjaVkg
XGejxmfJpzVXjgfZVSf7TMERQY0//3RLhZuB4YhvmG7BrNmz74tHpVYa0BrBX/V5
FuhV8BMChvtmYmatp2Fzc6Hog0pQb1QG0SJnU+A+917ECo8rJeURXiRiT3KKlvCC
Q/Kkl9RIqRVpYYrtZRIp6ybPyZkbpSPINg0si3udd2/UqLs8Z+SlmYDpiBnaPn0a
2hAI7WNWwUB2lf9NTx4nbVZl91xRkHzc83xEmcWKgjRHLVbjU1Sk23CUKLC0txWJ
WY1+P3L5mxFsGQXrUBJNYJA2aMvc4uTwTuix4ejqkXHO+Y6yUhZv1I8YT2UKMXAL
i1h1I49Roq1W3NQYRWJpMm5vmanDvcosrCLBZMECa2y9MZJpZ3tySUiPOA4cpie0
aEOEdcRboaFByD5k/7oc+njspxgh8baHIoebfAbUGSYbtCh8HEa2rDD5xMObkMn/
sbZELRjTYLzAetcaMFatThStjFXv6If+ECPmg8KBP9jEVfgPcobBwnio8A1k9o9o
kiVt3sn1U8BlTE/FfRkp6APBOQJ23xVHp1+Pybw00ymEPlb2pzVr95nesg2VPBm6
JTKCv0vyDFlU7ebq0w8AKllYLHtU62OgNF2ZvN/ETVc1w13ZrHpkHTs/qwG1reS8
FeVXuRpcU+f1E3FA+oSfRnvc4X+8s+qpRFXjvGxv80CIIPTO4nwgrfdJZm1YZum6
g+zeWmcT9sr0wNEwCECSIjMEFsW8p7l+Y+aX3d3U20YzX2E6bbwxg+EnImTOQpsE
rjpuwTrVsOyQl7DPCTNpyyNAYodmCUI1Z9RCu9/4255MpH+uwvktmhouLQu6BSt/
+9lj2MeaSGEx8BkznfxsEWy7r/wILQ7ut2+2Jsno2nrrsZSSsxzuNECIGD5WJ/9T
cmIaHOdntwT69ptAPHz+ZdiK3R78g1AM/oQSFauS9U22Ep+jMXBBHf3S9d21XTNm
3bA+/6NwLS6mdCVqY93RHu7hTIUwdjEQWKuTob4RS1Nz5CT9n2KfDcCsuvApKQRd
rt6/LmBnt17EevAYb3TUTRcST9ZmEOAqKNZ8hdJZSfNnZRBo7P/IeajCso+NSzkK
3L4P7VAs0BtISuG2CFQ2YP2/LFHGD3/GQ2PeBF2F4gJOWPIDOGBMy1jjdP3kqCjO
DkfO68Q2bw0vfa/K6CpscjmpRdtiodOrRe8oCaTDl5Ju2Mhib0/3GrQaU/fnfYCQ
MqHQ31Iq9crLZKDdA3GRVJtY7J+LGXV4GmBPoqSrlyypxyICIuD97LNyDb8gTq+f
Ra+48cc4w2DsqIWOusGniTbIEnza8zi6kVNfenIshwG491iw1bKqux0nJWWN39jU
O63jowDDhc7zhmfsDy1FvUcMr7FTuEVJEv/5vwtkx8uWMi118q2G8+QaymKu4YrI
wztkQw3RQCWryGBYxJb4ruf6SrtRp3DhhCkVMMungfs/5X+/LdtO0WhaiXActWvK
vdbLlgcNByHDkMJK/i9VRBIP5gKInXfERGwIiqoqaw0phvHu96nAxXdYfKWwr7M+
hvegDXBNxTrirqpu82dycxqR5AWadnZ0sv9e/HoJX+gaRglaqjWRl4ZmWF0mlJFk
GnH9Aub9Yyz47hC8zk02egIPCltodgmaQUALzGgIadARTpKz4fRB+Atq1MQsFILm
EnvHObtTW4zM5AuJLaV5ygn+mq1doj5jAQSeDIDbqLA+PYOjaGqOsIsuK90bgaLG
P0hXt2y5tVAIDqDCYX+OJ9Jy4vREPfbzlIGZJHfoocQ9oB/RvSXgSEH6PcZYlSkh
/Jc7b3Q+Np3aaKQM/yFBez2ZFydCw2OtCWTaXMFOt5T51p5V85QZl5lN7OCNP7Db
gVUNx5OvdlimHHshKyyVaMBEfWHtD4JJvI0CTgmo17u/IyI6N223vrJUpBfc8mJ8
4WZnaAvUnNVPf7AiXVOI0Y69qWtq5VbrRLdg220kynB+eK9pwXUpqYroEfag49p0
xE/kKp+VSK7k9fucl4IB+IMzrSHQdAAAQRL7mT5gUt6cbI6ZirJ2fShs4DNh1vpw
vVc7rHSjeRmmBeqMwnou8zpFzGCCRTCyZGZvyQvF/Oh3kHRf3c3eL44buhxYF/tS
TZv6Y7F2Ii+o/qxWqgOv3u6Ea191QzCm3rS5mM75B7zx/st7xl2dxuc8tEnuI93X
5VisHpw5xR9BJv8AdyZCQ18QHz9Ix99j+eQfgbbAVFI5YUY0g9z4bVz+SWgDBCud
KLBbCgQdvadzbPr7QvDlaw9VcrovGY+cK+9BwWUyEXlV+HaldaMyiqAoEcqAR1Wz
CR8qR2X1/cWf4rkSaeEetdA6cgUE1qlBq414VrvKElA32LjIsmXICweOq1zna2Nx
n9VejlMwrsAmF0b41po5TxqM7281mwrtVyANydbNotS7j8y+VXL73bXD9MizplzG
EfFZ13+4SevorcD4k9lNGHjoiuzX6+A4LIZxnK5Qtxv0d0XBR4ivWvfD6NaC0x7f
A0hnTg+xn6QYzGjelCHdDPq/m8ofEsRf/Z73kL4eRZqqhYwmLaCx/zXmiwWlKUSO
ItStrVgH9vpx+glwcbs+6cQXx1vNDsoRyLURZ1gFC2D5TKxn8zT7h9kDWkfsqbPO
p+xEXIDoHkfW15LFgYgRYLmyEakAVGoh7LnlprZGeoLHIiNCmeTRJ6ERTi6htBFY
DA7gaveIIKlABp/ITEkEflP74VGOX3t6fH6eVtXZNUq2iMqD+APhR4wY+XmGx359
G8eGAGNgDsWqF9IgyjWZmBZPuqcLco8a1fDdnVZYVjEvsNlyxwtNn2f+YxpE0Snz
4BwokWTPPsLvPloG423rNZ6P+sAGzlVfojDWp6rcBH399zQg2wgERWVmk1bp8Ffr
mZrh35mTSekdzyuL3ZhkvHBBScWIWpXyWFHmsuM+OkDUTsZzV4xs0vSq2YbzRSjJ
fY7wiqtVNE45TSbNsA2jpuk9b6vZysYIUljQwWf28ro3lDPI772uq0aK7vsimWCR
2hsHMnyWsmtH2Ym0tNegW8R10A9F31G6sIVp8JYlYYw8xQOKeCME0Ws8iDgZKst/
drvbm6kvyacroeJAlvCPO5mzAYFz9aF6eCC39mSX636rULLZ30JvCCvN9LlXoV2V
DAQ/jvD7SmxqwJ4tG135T1auBWQpQcgOAnLdJYTySUUJnDWESPIUnu7d9FlzGlxm
KXN+GXSHsS6oOaxfbNNrLWCkHkFNKqheIfVhNq2kTo38od9HGeaIsftewjpQ511x
iyzB71FCNxIyg42CqKOdgzjrSmfWghmu0Q8SwEYZ9qrT3DQ7YCoQEgMSLQDno7XA
OH8RW/DhHSYE6Cvs9hKWWmPNXxFYF7GgqICJ6m155WufBeD8ip28Ryu9z/r+Oas9
903c/JG/lNkASU6H7PBn10VJ1qIZBZPC5cMe9EJiVx5+3h8OmQm4Ixr1K5gOHMLh
kGXCQaFmrElvW1oanvzeWKz35lgJzgBfdyMEChpfDsM8G+Ng7Ji1vfLPQR6DreWo
CfyH8WQuM5DfO/L0aiFYbgxX4o2VtKyaT6B6Ywt5O/tDnlwebntk2sTHAfsigYOI
8AbTcO1CxzC+kCfBfrH6NzBo5HhoxShsN8jltA/IF3D1HKgyoysYXNjhM39PYMzG
+6SdTsib2Py0a2pci9nDwh0VzNuafIvmUET4Hovj/DnUFdh4lva5TPKzqH6bn79e
MAetu/+EaltvlLmpYT6MMQWPvQY5ytRoMC1EYL1XKFFdkXRWSszEkTxFWKRq7BSP
rnCkYebm60AW6PJuAebpUsFB25G0m9Vabo1APpQIMoeyRmRv76pnt4mYwfqKtD1D
78IY70s/zJJynuaxQlsF1FaAtSMpaxI6CZMOoBMtzc/w2fKn98ZfzStpH/7M3n33
wTJsUp2fk+yuPb1VeLbEN1xMtOA9BijhelqJvH518sjAQtYKfbmd6EJ0BNYQE6aS
nH1iHF4DjRc7RRi44EyNx9xFTEL7fM7Aw2tdTTNcUVCHMHPYqfbcsQOllYh2zilF
MZnnPMzy3NNKCm26gIPtsC51hFP9xYGkt8PyU0rQvzifHSuaS2mVWeY0Pqe1DEjd
9SIBoxn/w6DfEA5C+ley73M9IJAxN+0QcS06vGliUw6H+cdjzspA3PJMCtUcZz/T
ZlMpCNFtWn/k73uCJuh1U0GF7bRYGZliaGD4nVA3kBECdFOq2CQZ8KUbWvSM6Htz
TxHlEHNoZMCzvVQoqBPKopZX36cw/oDQvcdBCSIu90YN/17Wh+HEsVH3pE3+tvuk
jMCKoFla06JjxI6lCtBo/C2cw7zBXz/5PzG4+8emz6KqVEuTBMh0O46bwTOVXTrJ
Gxk9XuSeZ5UFMuaAIzoQ1QfFEcpOPPy0g6FAz0DMfZQArBDDKVyFTJ1yyUUNAo94
jVqxx7VRR5RFsVWyX/0W34lUPWHt30k//7BwGzfgIEyZQoXTOFKxfATzt14dOpZj
SyJlInjt6Ba7rllOz5xWh4uIu/oBASbp3+zH37Ga2R3iEbILiCTgc879kbsfT0Gt
XL7wJDX+AebzASC2MeAGMgtnxDPzapQY5rMyDEsEqRCUkpiwgmLQwV79CxxDjufl
d80h/YJuIfLvOZjp48cOPlC2kdXqvnws+2gLIxexzFnjg7dRKsF9Gq6aSYZ/1J/T
jS+aF910Bh9t4fehx21auj22an1ioKoCPJnmizfls0xvRoXEI97HLgsVPBFufl7Z
F+JMinlamLyQW5UWj/dWZWozu+GyA39w3CMlAuHAUX7fRtvG0XUsYFjd+PqOKXq4
AZxQVbgBW9lIuppzLu2VAVy7z9VeCwSTjV7lknfJFM1sqtYT6wP/0Tplxzug5DOw
vGPS2Yiqj3DhUFsqy9fPWB0D1N246Kn24GPIldgwvo+9m8JLPZ+RdmpnNTahHEZh
3Y4cHY7QVNFnv+hdHhyfssjKRiXsgwkpOcMcHE9M5PpoIX9JWMbnh7mOxV6abP3K
H+DN8As/vK03+IZiQ0L4P5BxV0nJcG0k8/VkbhhKi8292YLZF7o78grj/H/nE4kr
GsseoWzkNFUFOQB3ysE2C8GvOGo4ycXA+gqruXhVkvdSqHjj30AbBYnirtWdgwcL
2YFV7+S6Rfxoyy2vgGpDk0CWMcKY1jdYB/9wOwxUDDJTFYIx2Sdhh0uaoaARHgie
P2hJg0HyHWC4chkbKbjz37hB+UnCZWupotOGc0BLDq2jjoC2rlEB9z4jF6cU5M9k
1ZGrYamoyjMVZWJL8uokR1PIvCYbfouXVUNIKSsA0KaNpHNlwl8kgp52X5uHxQ+4
nSI+4Q6COHM6tDmfboWTXB8t+GJ//VayMYiKPtSr6A4jZhQ9MRpE9UOGHByiqjnZ
jzXgoXylQ40sDWqh7ZfXS/rZHm6sLq/SByEbKUU9exP7USsdjAObui2d+kb0WahX
BKxWf74qAO66bPTpdSJhpRN90vfki17/BB0LxMxUGvIXp2NIg0nxjsvVWtl6XCsI
oGa/xl/u9NN6MyVDymcEv7GH0a/PAxGrnJnkNE/sZED789shKNIRhhGM3q1xpm4a
e/KgHSMlr8guvw4YZsCU8OVCng5yGQOXEClSdq02Hrimm91CYfl1M0cfGm/IvYFn
ON99fRpoI7HerKKs0icN0/B/RzXAGOgUuhGbNXUDqIoXrVNJsAn2MmFUE5LzRWDa
U4YUUUXpR0lM/yE9+L3m3BhTQD3d7BE7916HysNgU4n5UMHrj4Vbz3BbLDiLeBlv
UAyyqCl7cVuwg8EulC9NRvMf2DqaUc/eYi8c2Jv0JMzA8p/4hK7oxi/5c/EoRj7a
7NA/GhITuyyAjxYNvGdVaaA2Xbi4de2nYOTzeSvwdD1Igme6x327/aaZq2DuDW1m
t/MyfSaHxhH79AGXFozAFQHoD73mNJAgobZyf6U6JrcT7tswAER5z55ApbYOwHT2
T+K/ePl2b67OdGYwyhucgs78rXcrEDF+I/z0jnHAAwxbNYLzxiuz20VvMCWyXxNs
mGgWE5n0rImaZ/+O0uaD18tx0+qzaU7vefJdpLc3WGiJNu2Q/yhOAKc3uLXTtoGK
A/+x2Rv+YUUQhufBvqGARLvH8Jm02Ti0pUkObS+Rh8HpYmvlkYgwfNXjmLhj3eKi
MJ3WOJn7+uz9SmE1j9qPMu4YKL2hinJYCVMSt7wSejzEE1wbIg+le4HHOMpliL+P
hrthXbxkjlsLppSWt31aoaHTcfRW/NWQkDjLi5/O9EcvqCDmA87d+zHBDC8wjfz1
ywFZU7y2vulfBUQEUWnDbV/sSi92VK29eUyNaSPK+8hYHrGe3XUJkBXsJlKzkLUz
6sx4r4LtXm6H5RZ1/AwN1cB+zWcB4KhrFRdHVD1/6Kuqw89vNduBBpVv3/9NxZjR
TTIsYZkKiDQJZF/rqtLmctsgvWU+SqEue2OtupGSkOD2lJvvEyZaXFo3O0UEFwAf
jQ6EwbAv/aslod/jupGQIBWFDMWK+OKlg0k5v1vvNw99k7nJMwm/Dolr68mdI5yK
V6dqNg7sS3ptY/DVBgbOepEcl4wn8mh0YIpCPlDGQKtWHTtGkvEC1Dlmt4ecKj71
YMTa7MPVz5MNXDW1JzRWLIurTx53yoZblS2cP1sPx5t3DlSZ9UDT6X+o/LTilwUF
uqJoFdMNxEVYmVZb2WcQnpOOQurTNlIoX7sv+4qPvtQcL9fm/geWP8QorCTdsKuL
TTMCz4tcjF5MB7lYdLloNSznKeQM9TE9LA5Pfrf73B/Db4PWB9WYOFP/2lzIv7/d
mmT8gOHidh/ADbANPCEqAXMjVro/5CJA9UEeamtUixGMSjLZobhfU6miHxkhQmCQ
o/gA1YpRihfTpO+3WZtt1ouLqN7arl+RlqEGMg81yp/BiUKpywVf3VTgMh3QPsvS
xeLg4j7ttfL8k8P539mxF3kwlk77l97z5dL9EIsWiw0rJVbCpAtDVlnwFU+SBeC+
xAlqBztNNqfBVGWDhft4AUZjpTUGqypCRzhzsTVfwqAjV6LS03e2eC33DKOD6ujz
NPpkBbo8/v59CDI/ngIubZFxrmK8MsfjhoEWYqGnTdW9e2+QmKguL+ss2Caiu95H
As1d5/mZw9aeoSvOjroXWhua8a/NmX8djAbHZc7ZjRkK76NwnMZfnWu+hwoZnxfq
0vXobMJUiaV5CqmJ3n1WFwc3pdZQaU/U/pF7lsRv0fW+tytG3muPopC3huD769nc
HypHQNX9eMfEIKOw/99258aTQEWy5HNvsP6Qe7tBYrQvw13+GYycj2uXMJS+b8Xs
wZHJYS/Fqi2hTzuV2FdH3JpD8NQAUJPs0zZBXJWeYtuK0EfC/u/L4E8ipd/iFZlT
t7a6IzObuUKGds1QyKmshnq6XNS5uiI+TX+YTPbr0/MyJHe+5HbpCzVw0qeHSdJi
JM2b5SLuc/4XkJgPSXiF1IUl+t7hZM1OboNjCxXXL39ESDxzlglBm9ulpbCW/H0z
YkZTeB4DP5e9zEYN+o0HiLcKkZQri/YgFEM+d7nDuKJL26lNZ0pOvjzFdwvt1jzT
4uDSOXXSGZXMDQkHXGsZzs7KGTS9xVSGqGaaCvYDspyQH8tyvMEj2V1zhs4OlmRA
M5k2BfF6+VZG9jBAvkirh5ikxWwTKPOo8ej4v9sxggfV+Lf8rT9W51WNqWO5+CQs
BexWwiHq9/Xq7N9YmO4FD+lU3Yz42N9cuXXNG2nkws1ZEBN9kT7eK/r2bckDyH9Z
DcRcpCRgtSBPXoTgYZKZSj3vU3yYHlkn+B0pwrxLcFBBVVfm5mtmySmQw3SjjRmq
rr1HYLUeQZH3ZBn2B2uFRL3tRNKODZ54Uda9VgW/q2fFRGYbhBti0VXNGEMImfAL
NubyBxFl5xQLcOYF8vVrteIOAfyBNT3QQHB54vOMQ+hLWacIFqvZeD/uhWR+iKwj
/lTHEs4TZAYB8NFBHiRv8ZalBJwBdKuN6XJpvLrU1/S0pYxXrrJPVlBpVXsqrRH5
gntkm/S9xyF3AFYFSLXJiqWlMxQ3c1aAcYTPWFcD8LCiiNsmoGvJKPmXO690/XE/
j4QLKfWIGa1VXs8eIcz7it/EGtWL/LSCYn4pQZORnuLC+cRlFEzp9ltnA5RrJkN/
ekg5Ss3RdGEumLkag8fzTJkCDUI/utB85flA7R5x3bsY3FTW9H9ise7wYLHsZVpe
RRfntspr4J5wfkn2iQbTbx5mhanMEa83F5FMYQCGlPJWqoHNtRPJYmd8MYYsuus8
UoDAhByo9edo3sMzZuNexvgH2/qEujfCP2W33fNJf6ZyozPqh0M957jVGy1nJNG1
8zlbyCRrjjLzlBPXh1G/vz7Mia+bGFBJPSMN6jNgwwqShaf8NVTnupuwBAVImaB5
5Po/8E0S0Os1YQaXzoYWdYnUW8BC4Osgv69mTm0dOXggkCLL4M4/hDMq49CyzaCu
+z5kHAbH0XM5Unq6ZhxkaGCPlJ2a5TvEsyvNrhC4m3qauyXcRXFR1nTpXTInAAOz
65B2ap9IN0CC4HAfNhMqbwqchTF6GB/KUhA/YGA22zgW9D/CtoG1xJfHFhbsPW82
JzXcdFLu4EpQALrd7avh2sQ+S5gDwPX3WcGYznMN2ZAJBSWAQcGA2g3KLGxkrHQj
Uz5wRDZqCZ8iHJtKVXxJINjbH5mTkfvcp9FbA6yIuZqugz9LH+OFewOeHHRsJgfy
atbrYqKnhoRgRo6uPdsoBN4+EQLeQqRND8KdWUd0eumO+fiUWut/cOrGemDURBEL
nAmX509UcTfZNineSeLUGhAAo5qvLykYH13kgXP6vhH3a0bZHZnvpycoeNg4KX8w
o4R6d/Z+4JYpnsN4O0lN6kIkmnInmjpb6/gMwRKQLpduKONdaRVg8gtUakyVWCfc
P6OlAH384RWtzCvpFNtNRJAWNIXT0zPjOHz6GgGdL3UtDT6yPwHVahri+hTANcgS
t6M34RE+ZyIyez8FJ/T+Pl3bpMqmYOlc/wVtgb77rLt7TkjLLeIbrWuV5cIqKTw1
09Ug4r4CrURU4kErFOaTzRc5UxliB/oIPye3ywU2DxL2+1lNyS77jNW1UM1k5pAA
7wXRAad2q3KzR51DH/pSqlsg/XEkASmn9KaOdcBsA26qM40+Om1kIS5k7aBV6h2e
zosLu9t1v10XhH9XTbENcat5Rm94+a/rD9wxQg1BJWJhwrTytNiSI2e5tIB/bH+m
TdZKmIK5SG/x9PN2xOmqtSN0hHp66mZzBSx44vQkBlRgk8hN9NHRrTZg0EJzplU7
dfIMXPZg11X4bq6wVR/e4stzhCNKbPT4IjStpPeucp1ys8/f29NJr6cgfewK32u2
JdsYD+beGm9lw4x268anfHVg3XGvV0T8pAJQI1nwAN8z1lpgk6W8gGgcShJmd8O6
OWjokIy8Hlp9vWhwLa+etxHbgeZt7s12d3xStDrNdQSWO9tpX/fZhyOQ8vP9wmUt
xY6dXaIVMTUQp9kiQ1IO818CTDt+QJB3L+1V3yvn0OdyuYs5kEXPcXbWaOaJKoxd
7GwNpYS7C0xG2iVDyUrq7jnNF4JFGpPpi5tfIbb3wUPO3QLsx/dNr/bsGCYEybat
kRT7UOGtS4H+xhDWEdB6fyBvwCtlbN4+MYN+HHHiLFhNNwo80SPdqnxoDFg2T9Qn
GG7RprHzm8Bk5ef16kN+s9T7l+PMJXVHG8U8SPjOqY/M7NpQSDpqNSnwMA/xAZ/U
1vCM4j2T5UTeJc63DRgTUwieR5Pyqb0x17AHee+UzDEJHfzUSxNHCs1YIz09HcGa
BMYziwBTEta7upwqSQ2PddRfZZv1GZaHBJPjRbgamSDXqfzdTMALbloan74JyUk0
tTHEwIzRYMpr0MoOzUJDJXAKkinV36JAOSumV6Ockvh8RB0GnCYLMg8HPCvoBKiH
Kvm002FvhhgMYknNXXRn7D4FUH0ZYnR4rl1sR+iEFpm0ZdoKLvVq5jgGKnqhTyi/
n8NwPLt0Si2ctg7llJtwkTMLkDDbKuL5enAPZYHNyZOY4ptzuxaKK2VwVNKAjIv9
UpAJbxL9OU3jvuow6DkcL6Roa7cS6PQsk3ElpPZdvmIRbQRDHoOhivcaFwp1JL3+
eE6107ZwYpzahS7HuXiDP2kxF5KlCIBEwn+69bWQDZgdU9Nb52CuR92yRj5RB6/E
oCSj9km6u4AQSBOr+6/Ur9gWiUv1gofopzM5HGI0CZIhzmoqi1+T5uxOextd1Mq5
nTGTxQ4kBgRoiqmkc4YyuiOBcADEgc+MAZ8Al7V8h0tI7t+uyIuP47knqnTHUKeR
OWWPXsuEOLVNRS0/9XHmqDZTw/KbxfZ5BepZiTLYbLxmhw+KYgN3C2rCFgGH3MW9
i/gZlVz0ZfI+eiMZLRd16VDP6xjEnceii6pRhfvN8rRnD0wpZmkKC2/byVJs7U0g
r79hSZBwypNglLiS8+NLP/Sur+03IgsWKBBms4wuUpakgzgVkJ6exU01zTnsxcSy
jjdHrZM3oTKlwAO/VIuj133p/UlBRA87SeuqGDW0aFRoQDGZMtQ5nsQybpzv6Vuy
ONWgNbKCcRniJ8q9ElDD8u/8k89owjO4lfQP/IEpTieZldkoTHzBusN6+ql+8TNe
ZZRxjr8U563tPWgO4IYGkp/RSnCQxSGZfxplR5uFC9S+hkYP6VT7sFW+L8kIPmV2
efVVMD38GpXHBEsr/oMAwvje0edGhauqWOZF1tiTfw1NIqAaVaAAUTxmiTaFCNxb
hY1pfIVnH5Mkxrr3Hb4iLh8LqZCdjCCPeSgdPcBXUwE5/cjrXjhFdPrGqqantvXS
Abgo9uwYkaxQ9DiXshQS7bW/W48fE/BDX4bSdKjeD3Ol5suJrRgxRsXD0xscqvXT
CaLlZru/0Ex1ZDchiTe9v7jlBNdMw1tS2qWYHJFixhZObmGJLaAopdjKX/TnNb5T
RQi8duS0qR/59jioiYODAUp3eDxW4qe8+yenyKfPr55A0L6EdQxNEFee7bq69FPx
BrXkX52lxWHwidkNVj54Wjs6kA9+uHrRI2wATqKX95zyXrhaBtIaGHaCcg7wmvuF
I5vEAEGJuw1MMpoPYM7+sr8aeVCIYKlsy3sNAQF4A83gy/RN2aM5xI2M9j5CmNT9
pI9GbWOq439f58zlSx15umDRv1JGFvsLLhOrxoHApsXA1e5aUYoRr2HamESCHWaU
3MiWErt2T0m5H0kWwoSSz/Mxbpb0wPKji2qCyROpwYmCfoNQQHSVzDBvXw2dgfrP
GXinRHxKVMXxlWCkDnZSDN1/wa33GPpxjjAxxH/1b4cwCf93i84zYLuSi3+pDH5/
efOQE/3TqT6MSZIWrvYbajxZs+lm/hoKBCBR3eSIF04V3bTK35/LqdHc2XDOKOx5
hO7r3KtIRwaVxHPDYBoW1LxCAGt1IFiP41Izkidkl1BeRe3bkeLTSDOJUQ8JQZSm
4C3SYAsUQIp+6RWOsfdzbneuH5EJI8PyPXOJ1XNdb5RpUMy8hn6daAW9mzCtCvwR
YWijFzOxLyzy+hlt13pUw8T78Qb7ToLkf4lDl+zekkdR6vw4wkUXgHi3f2OjHF1Z
fPotQD98ITTZbROSKsmFvcKsfGUcvrfTz3sim0MaXwrOm6143Otr9zY3YoJp7XDv
r3b0p2+uYhMJ7NdWUxLNajBEkRYdbmzWHfWW1iMgQ1wLugmDIN1xJWGqguJS0TsW
OukB/VjviiQtB8hc7LmPT1mRZsxiGzzDxc4vgc9vr3cfy8fsrEbZa6u2zwch7nf5
74BOqh/FVMIBakXjEt2WgSyttZRo/L1ai7RMLItVOKEmk2hJjIzNEJgCokMWAOYo
38E8TcfeStaEq95PhStbiP375FSRbGE60EnMrSR8ztdKJtR7Hf8kYgREzcwax0tW
6kdupPDJcHowEdPySlEH/ce0Y6Bajr2bQcfA/BViywmqo2QlbUAqpV+drQJr1OkG
A+Fi9wF8wxAtv6kVp0q7e8DoZHV7ovv9URV4URLxhPk0JSPzR+nibhkL9cVtZV+S
eN6avUX1U2ix/ju+u8nqWvYlJwUGn0rdV/feGlbFmb4fgD2SoWECbyGD5pWSyEPe
rxvwFevWFoNVKwYcDixV1SM5KclJEAKDcXGE/nD9GzWm/09/kW030VJp2BGyhRe2
XtUY2E0VeehVH1fHvjF/4Nc37HOKpQGvX7qCL74VAV2fZ5D88GIg+eGad2Mldkgs
rxtln52RTVTjl4eEfkIHLTMy27KnKun+JDhpFK1EFk3YWlcppDDpFwSi/rb/ICY+
oZOVEPO69ZQN7nJsHsPs1tcd5/XUSUkF1rZP5/zzeY8d0kyTmFzIaA0zUbipSwtj
uraHopaTfDlC6eWzEPtOlbpWQ6GW2wSYIOE4ssMi4CiXnAVdWgqlH3cMyi4cqyiM
z4VgKrUBExf5vlAMbbYVClw+pg3XjXfB1LqprSRQ5/frRBJerelCoISHaFhVMSkf
u5b6NX0WsqIVsNCF5guV4yg3YWceiTTwtsC5Cby6m6Kj4y9qyOltkYp+3jtFQEnY
P5tMR0eyKIUh9mpOryhR83MSEJrK0FjfifJWixeZ0L5TW8SEzhbor9ubZaTGw7Qk
0QijEdUtB7oGcIuLoCHkPaneYvpetYI0a3OAGW9BvRhGI1yiefRaGBG1hdlY8/ny
iJfrXftKmXz1zBGf71IkUWodzsKe/2wPvY3tZdadAOGSVFiBrUYjG2NOiJM0wtsE
JRzJNypYqIjFHYdhcp+KCDD6TkeRbIXE7fw8pWBgiFePDAjKMwDtmXo2/fAeZ2KQ
+bbjhpEJgWxsNib3ViJ7gXx7ZZSTjkmPD98PDSnKBn1LPrNPLl0XruLApbKkjKJ5
vMVZajFbsi3l3p9TkAJLOMYTb22kd/NbB7rYkvhr+aGuQSyyZ/gXl+V+KYrDsdlE
DwAmp3t/2CensWkkIdd0aUYn+wxWtbhvt0LvHysYTeYryz74LNjn80NDldTBbhzb
e1UnKKC0vSdlIvDbl2qBIFRVmEaKmSJVMLbtVZGcslX0VTI62tT2/Y31fsGKFY85
fcrOYVCSaZQwUG4ZGjR498BO0S6Ih9lN39PSYU3x1s2pJ6PWvW1Kv6uRVORlMiY3
yNyemWINAoeCO3a/4uR/DPPgrXalw4568roIWIWpJ8HIJzo7l1BGghM+pL0E+McJ
br8LHqSJ38/SJLkDV28g0g+iiDz4eau+7TBKKXMBN0e1AuCJIzSvRhHJfo8C7I+V
uupXdnWYS9oiTCUBcK72NDhSSxAobQjArmZ3GPiPNRMxhyfKeIc66/BhbaiySwG6
F8KZQHRlVtinJlyf2nmJ+N11P1L8aJ3JO8/Kk3cWmFrXL9pX/35Z+TH9ZyyyObp8
307bV2f10RhFGys7PYY6qU/oHNRdqqT7puiAa7qLuLw1i5lqHMFTD2rLvTXF32ER
oP8qXlIGpPY2HLTL84d8cwaRN8ZosIv1qGxjnip3JQYdbDHDA0tL/LzswywTYHHU
FnKbXu+fORgH+yXoilXQSD4y+km3G+31//XENuw4yRQpAOU7OMdWFSRjKSJEJFnC
6CFoUpprjCfcJVI/c/vwhX06PZh6imkJJcusuU8LWxQ4z+tNefjMzQkgTbP/uNeL
rLT8ehOrC9PnDT9EdBmcg6Y/FQvLDySobxQH5RKIe4/uKqXcLfnY+Ca9ZCXbrgTg
1HDsj0dFz219I5fhGE6S6VJHJFh59cbUapqPAOirgq0i4Cv35jqtZB+Ks6moKI/Z
h9KD/jr5IKhdzURuBvnV6R7Y8szh8ynnOGqO5fdd0ChV+uE675I0d9QaN5jYwQvL
Ue91sIC6ACXAZQctD2y4Jh6K476/jV6b1+HVe5r7Gq9gO1U041/QrGV3/3o5Ldkd
a/GoZjl1+ND3/tu9lNyhqYlWSOq350JngnCkopseuCWpxmRsBn7hMeaI32ywa0x3
s2+xWVQOhBWT86aGBovzlV3EzQOCI0LiWsOmWF3JUyew//dLEH9gHKPojY+vYQO6
jDdoBzsAtx4aUFAl6oL7Brs4LvSd1obxILv53/v7/vSuoH7OFYq7NSS6VfOp4WJa
DEG8rNDDdmOahGzRRP3EOk5xRO2ZrdItAnEV2In229ta6yXojPpGwadjSIqHGn0U
aAViiRAsdQDkfm526rgJ8xudTs9liVGSWvrONR4vESeDLYg62TkNHV33ZnjrFSwR
rGak8nMrdLREMfZsli14zpFjl+6sIaND0wgCoH6i4SQUPI+m5DgbJfCIDE6HeWbb
DG9+Qrs1VrUD1W+tHtFrqsHCTTkir90UJMGRDMHX1h/8shlzRNIjM4W8fUpv+afo
ypMOxLZGGH3xd2WMVPB+EBLoqyXhMq/NF07pBySJu7d+mYtgkiaGRMYJA39jMJxC
fWDzhWocc8tsUABt0UgxD/JZOS5Sm4TrWze26hx2k6O1xwqiAO7wLfUbrfIRS4FA
Juo3Urnbn5SK+Z2N9PfS2VgIR+pvVDRL2Otk68ihY8OT2lOA+31OiZ0Ony1QDA3a
eyG7hzJo/SUMbhU0wByESZTaVWPKB/cekLpvS9K76JVCwRUEJG166PzRw6UG8zeD
NCm+x+Zpg4KCIhdALWyXIOXpTWgkW2hy677ROkjX5C44TSHlb94Q3BN/rXMzewlm
dG6X3gLKvRcY6a5ZsMBiIQRVSjxUK78mEvMWa4wdS3hSCgLxllMWKufnPJ5Gr0Bd
R/V6s35Py9vab3vaCXXozHMIXIW5x6r/lbVu29glFgDxrBuzIDr9PVG4eNaLMpy4
8rjvkW55mEvv2X8yx90KqH9WUZYZ4cD6oQpXOgiChYH8TZ5faIK4oCLXYVjhsKpu
+x6EQCQStzpTJXjo3oKQf43VZdAdj5s1n2sk2ikmXpXThmfKQQir+dks9ifqs1pR
DroXGczDQJUiR61vhqZv1KlPjxLdI3IHL65MrU8sSS2aKbS6QRiiWTzI0PCz5gJX
I1bMVnczqzttPsMxW9F9XnwIahNsI8aa0vRnHUVa9z4cNtU1sbGrnY/vBLH7tn4L
ywrZ1f4aXzPIHD9vQcunv6hWUE4MB07eBKW7m2JabxWMloHEv+JWBK9dlTuPmtnu
9OWYGbFtldA+gDhunLjY1Se9JvnnLNo4z/yxMps/YsPoDnOGzyiFK+5ZzdtV32aH
cxo7FFwWHpTiW4wsR6jLagMF82jGMU3eX55ZtP8jx2I68ewzeW22/7x9OhMkdN8f
ynE0ZEEf7xqQp6z0nWDVQu+JTiiBsbRPB/pXEGUJAjN596ie3TGhovC01NciTZgr
AJpmn1rV7A1dPUSBFLzeBqaEDkZthwlBmXAkUVZl2udm3oeQZNRD0VQDBxg1kOaA
QbCZzS4VkQenU9x5sLnx0bWtKHo3Xkj3ImqxqSLhXkUpgs7lItfmzPSs2kgmXhHG
h/ZjrigpJLaTIIRGFWxBEv6mnUGYMhcoi6F2dnI3A35QIKKvjAiey2WfyKRCI29S
PFMPkk0CVcNoEDSKjqzDk5DCVeAdA7XS0HPrMAxGBfeXtl2J2GV5vAkbwJh/0Gc8
CxDEbSzsXFaHDN3OXX0NZO3tKE8i95OzoqQFsqCRZTisMySnwbtvtL1ApKs9QIh8
xKxKHxvjV/iXsocEnK/2p7pNj6VMihcmet5sPQ1D+HoOVSvdZP3O1kZoZ7Ims/zf
o3lFPSfxg53b8bLfhl6Ri0ZiwFeNvoByNLScBUc3pb9cHrGwS6JA8/qvtMMDFpCL
szpjD81UexJcCvcZ3khnHzkPAMwJBiLhLMiPZlQRP+vBfodEEls9BnQO0/KFev2u
yvszIDkFtzk5VMoI0Us4mqcGl7AcCpF4qcBdZik56zRvzKej0zDBJgUjWBw8dpHl
oNdnhTjzTkSuvzTGDOeizY7dNEGcuIM+xiV9opWjzNVTfEQicSl+Q3d6T1afo51f
8iqkrr4dQ0bxQkyQ9cQ7UJ3F8dXMm9U3yxVfrNoN7Lnf2mxQtYZZ9Ucy+9QjUecM
idIf8vAf2tInzNLiiHpB/NgYiMu/zx/K+LakSfBsF/Ljb7LTWG2gNwCF/gEpLsBn
da/YsfWcXG8oVBiHQWFa+4Lcrlcujp3hbB7yRCZ0cAEKBVV+1kbxrSdJp7QSkOcw
PHpzmkRsWxNG6eu/Glx5BHByXVd9fegsyoIKQ4J07WRpFPSAvvjijn1M5G5KJ5Hu
0bjTNbGazLdzli9hp5BufPZgyrqidmtqDQV9JcKfq29zGOmoLzDeEb68r75bL3cg
VooOi5k5bZXkmkKGZaITjyEoPcg1w25aYQwwhYOZSR38+1n6ETUeOLx0dLpufJ12
6+G/UywKGIJv2J42DugdkLI9sMzTOnY8q1Ngu1P2PZtPpmMJTsGmUII1c+gq1MiI
tM0QleIAU50TYaqglHciGyjp9dHTs2lXOR4JfnMP1DZ3FmNHBdLAo1rItUyxgY/7
gGFYobc5Tw4oFcVX637MoIrNQou6Gga0Lack5YZKZTIzX6XcJQ0yCNhFP764vNt2
pYcg9ok45d4rMCiXyIRDif+bsvfX0MrKLwgp11fiDfzoUdABkKsShPnThSgcUJWi
XHbtHXOxomaJWqeSu4XpcWcqe7190JtlPlAJdXpRbp8QcyrOCvYYeIDjF1sWM/H5
HNinWUai/ALzhWETtR+AVElCvJPLZ3XlU6PjlkV6Yq071+hdgXV3FsrQ/f2oz9yr
TyRSFyx9xe+wl2uAzqnIQtCMoA0XFer6H05itQc1SK9uCcVzjfBQ/UlsXGPi8ZJO
RZwDK06SBg5GT+CGn44cDTRH7eVMcnjNU5S8kfsCWedzNJw03H7U0Y3LctGsYqq0
oO/dcCkOIfD9onHKxGreRj+bwjK6l+z6bhzXWLQp51Vin0rnfHknGe+iAc/hc0Si
T+n25VQDgenwyy3ghWggMwUi5FXDrq5EvmIE9n3qZWgU1TGxW5qaSSkOhZARxDbD
25l+xAFihcVvSTLaxWUNFys8KPXz/jctWUGZuwvRuqvdxaq0UNvQcZ92Z0wqGFH1
BWo9Ef+FSeKWv3yi54a67GWYEHJaGOekL60pP18QyjNLmXbJ0LAZo405zcZsi9Cm
Kd50UdxnmORvAPDQ2UMwdviKm2DODIJpydX4zmJkweIgnwt+H59oyHwnubfi6Ih2
2ZgS3O2HKX+6fWIbS5rByr3Ll8Mdej3Q86o1BiZCK5qeKLPIcvrnXeoqdwvfOdMr
qxXNHxeLCoqVN4X3q2wveM4HoWeT43eJj8MB9m2pdKZNHTkwDuwOpSZOecnVvUM1
mMMKyGNq739WFAARpuTW90PC7O0ey1GRrF4GeVH6IadaLpUVwswGX94NAi1TkbJI
zESqBIZCFXCULSG2tCwqDLj6laqc5oadSSQJg6CJbOoG/J4dMsaBJ9HHEr8KpoGP
VpgbOz3Kimvg1gm8UImZ0TJfwfOsKoVFT+IAtjvtcMSj1Bnn33cu8OReicOZDEyz
QODuNcskRoYr3Ik/jii84RxRRkhY/RLuz1iKf4rQ7Zg/iWSYpXjIqqa9ze/8+mQV
F94oQgubI7KCAqZbxiR/jcHoKjisf6lvb7rBssSjog62soDa16nYUPqefxL+PZBh
9fs2WyfbDZU0+8MVF+LPK5CJDaCIXFNzT6y9668I0pQP7u9WfZ2cgHWLO7y7NW/T
XW2b8I5ndPjEllxlNnmWrO1JfSK/05Mg3zFNnFZE7rSEGPyS/WbXi7Yk/zScLmRJ
wzkgLkRD0OpobA/UVBoL+ki5XBHbHgpfV7deGutTkuxDsr12uzn9EaLxY7bmfW4J
AoQyit3vGQDZugsOu+PyAfaAwCBnPJqNdJGNVzUaL/GJL8cqlsMSPBzFE40gqZlD
Q/Nwzqgzveo+Mbrwva1YcHxjFuGmpnrG/UTDN+eM1w0VZIysFvw24agF8p99keQs
3deEWEw+ChGBRFj6p0TXzq9VZ/Fbe/F472+Ps2P5UFcS7+qSBVibLQNRm+mEgrmK
PPEF5eviX99UbBEXGR6IaQomJb+jJqp6euuIJ0FKQanhAU5fFoNAvYZZt1PZDRJm
qWc+CoU50sskoJ2NSqxlIXgY2DfyANoVp2hfS/nzppk=
//pragma protect end_data_block
//pragma protect digest_block
xt3Jkq2bA2bMX/Y4Ra+NHbbQopY=
//pragma protect end_digest_block
//pragma protect end_protected
