-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
sMV2aejFS2U2lmjffvS/4rfsbKkir9mZeHeRY7JUrCuMkbKpLR0LID8YrXINPcqx
AgW9waaBhlKfmu+RT6nERMlpAocPMW9SU+C11EibmiZyS20U7YLxtsiYy3cVHnfi
rAfYoFngaepfSC0nAlMih9JnVpdTou2c1cHLZJ4dQ33qfncWlXOspA==
--pragma protect end_key_block
--pragma protect digest_block
tqwIEXGv++P+9AxfLH5JmVmjVNU=
--pragma protect end_digest_block
--pragma protect data_block
hPt/xMl905URiuCavKWkor5uwgTEhQ8KGVxWL03MyNbGRNyjw79CfQB2+jy6jK50
UEEprHtIfbQeUCU14FrlaMjSmvwWv3cD47KUuhJrrfV2zTg2+7ypVH0N81eJ7SfX
koC0sLrqpoaisfwEdE/4S1fXk8YMGGfsPC5JcPaY9Y3KLvj2bLX07FFzNdTWgtZo
oeiBNlebO9K2dgZrub6wr4soIhfS3rjPqOPV0OuZaYtGoh79ozJvNyPPH+8F9IhJ
lFXdkurtOiVIe5Aexcm1a9U+NvNiF1MDmZHPfSF5Rorhx9/kP9uVx/lSpHu5JldR
OKXstq1hn6P3C3MsQ+LUw2eXWRzcjY6OlY7s3HaFiE9Bany+iKNUNSqrTnCA4E8F
JMfJq2bvBiSpv7YA/3y0tHWQ4Nd+VvZzlRY34krAHpSuZ7hn23tc2Y7lZZ82PEsW
Ez0zPj7FQ/s7u1IRTLTitLXHIwUkpmHggchTVV2XgL5iSRG/sHLGk0gx1wnQh1l+
RMc/kEP+DejBwTgS/XE/BxUgMliwHezavsxmbVRh7dbWc8DCqm+Wy10Sc4gKdz1I
ff3SPSxOnzQjLMoNM88EOUkz57YJ8VGE88RmrEE6CIh2MBJz3sfNARN9BLBRRDyn
1TwX0TwuP8df0G/5fRvtf5fRksUDoj5HtZsHmtQ7WQzTUMoS+qvxyDFMc5uEw6st
5dO1ngOIemowvqnoJvMmgrSvz9M17VSZCtvY4K3Tar7RbrWbgVVo46jJ/aB+2H53
hfrTWX32lyDEEw/pcnFaGZpMvinji8tafjMoPMiR+yuB+baFEtRbZ9CS4RBlAzFZ
fpg6B7Kclut9onydhZf1+gya8nbO4F/86ejCr0wAXdbqIhqVpFUata7x+29wCETb
kXEzgdIWU8tVW4iiEVVrtI7P/jcmjauPn+aeovo8m6IvOZ/ZTh302ijd4HlMlZf7
42vrX9RFN/AlZf4PPzeX6gj/5LXzhNGHTe+LEwZ6y5sUXa5XyJLfpcjpkfh21MAu
bov9lyV+U9gZpKt4g5Z6NB0N5uRYdM3MR0XKsRSWx6SG5QFq1hWjXYLBbzxrF0sQ
ENI9s/lG1Bwg0C9I08NxzHpbsO7tM9ff1RQ2JHiiNWwxclj8NV4ZeJcvPRMynr9q
+nP6mJKTyxJ5qTN6AGm9vUxW+JIhk4RZJoxwwnFG20hqt7yokW8NBitg4IVgp/bt
ELlQdOdYBlq19thY0+NYV6xiPjT91wN8yFQDtu8iSXH1by5nUPnalVslZtF1PqQl
Ieuo08Es2po1h1VsZHGNQc630D2UQaua4pKgftWcTMA9GlZGdbhQl97L2AaF1n3U
ykCr2VqD+aa33aRWNv10UEAwMyPtnkrVHdWvN8xrULQHe5XWXOL7lZYT+XXA/yBC
lXGgAL0vevsF93cL78E3TaM7IpYjd8St7PGqmF1ZxOb3URduPEMlwVxH0VgkfIP2
ftxr3IeX6TcJ6uckkNefFrhOeiU+kv/ZRp65VqBLVHaduGtOBxliWtQAeyuawVQc
tofd1LxKXa4hEr78suvw/Z5dxUhBvScFXo/TXBD7xWI8u+0CL9GMkOaXy+eEXSXW
2wXdEIntHY/kBA1aT2kUKTyapxfk1Wr/b2AazlZ0Nc1ZCTQtPS7jIfogUaIFKW2e
7U/hgH3pPwsigL325IYOb0jYfuVDztUKyoTLq2xh6Lamc4DDZ4hMNrP4m82xu+Vk
cjI+oHEnzHL7mueAITAnc/2lrFsOs+e0Qt6arLKDO0fP2NX1vxJOmDI8Dz8cfV3A
BqHgZUEQvKXx+8K9G668ptkElQ7k1RaHLmtTwyuYc7bwUvELLWcDdvWBQ81OKsqS
iifQPQkBABAvZtooAAI6fCa2qJXoHPLTd2hF5QuLQ31tmedi1I7yNXYZAH0KhWR6
qGuZ++qDe88tLGu4eGCWPU3oh3SdHI4LQxOiB05gphOzBVJ0MOoDoXePBdDsdyUD
ctK3bnXkQ5tcHkpJ1IfISWyWotAfuBQbhBRbUVkQ8UikXtk+STsDuZ41PiXuRFo1
xOyuuFqqSe+3xPkbnsj0d9dQZmaZ9lFPbZNQEg4FBJFtn6o5yjzLgmDlhWbK/+4y
s47iF2XMs7KqOOtKdvTWthtE92PBVH7GIChgZDjuPTt7fBuCqVc+PHxWCVRMwT4o
IDVF14gfUzHNloKJ5hTUEDUQ4BsBU24UfbvVHGKGTRvotU4tvUrgyd6uIVuJYgdS
JW3wU3EWzX7b2WpXT0MxY2DyfPMJC1kf7vRFkP5USocERwcl+hdGPLtvCTTQncqV
0UgTfqr5fxqpMpS7y0JL3nCn40oaSsat4QVz2uwTGknMfp9OQHJ2JR7cLEbNNRZ7
ffCcrxjjECtnp2ZK4MMPvEVvhIdb3Iq52ftmMQCKjvN+QWiTgnXPLkZQP/zppz/9
jBtg2Cu9ekpxw40PkvtEf+UPcKXgDa0JQVfpfZSt/UeWfmXBkrw8uoVH8xVM5j1Y
gCE7MTeeuVdtGdHJC4o436iY0Z5kw6YGxxqaEqxiE0NImJlP9s1cyQDJT159yNr3
pbDDMA+YRkd+ga9Pt0kg13RvbDNJF/4BuGeyDOOFWOiehBeC3OBjNCJUatPKHP3N
yhbftv6MDuM5KdkSFV0S0Lb5HVBY+hLtnH3sKS4Zc1D1+ZcOuYcXIH5/ksFojzB4
wPsnMhpbGs8EscpODupuoUeEAEcx7Uug7X9n+Slsk35SXdz4aUZ13cxakHYTtVJd
83qgg2TL0mAginNr5ehM16IGFpTModr4ajBBc83lwCwlvkAqcJEfEXMHDCpLmZDQ
s49ULiC1AtkfYs2mHbspnc2TRTmJObwAr6BkO91+wqQZwhahPfu5SudMkMpananO
oN14lnNCLI0IVVFPHGmFFNPwHjtgp51BdNA//mBJhvtKPPy8hOEFokFztlJUQf54
4ziU5fumXbbRbyCCAPz4rjSuYjrAAb36HLspP+w1WZTaN4OTiamWVZqHtfv8n+ma
KSK6FeMV4Q1uT7+N+3EvI04qw0vDe1lT/aT0HPw8l8uAh6ougnhqSNQdX/Q5yCzQ
zY9bzXOIyeeRoL+PH2/exoOjt0JzazKOMMpKEZUGrMcIbtMNWYufUOMAUZbaxPRt
IFaZMKCpr5tjq+tXYnkRkzQxRi4eyxTVYK5DR4e2sMyKEUDxrE2J2CBHGGHvDmY0
rYDMxK8BPgsr9aKw7AobZVZFmJ4sK/P8sGfQnMABvpwv+f6oLt+o5Vdk4vZ1AiDQ
RQJztpQfqF5D1h2771JqmAgAiDhBKcLdqDtM1vTbVLNWHGGcIhTu6KhqLrQFQsYc
9MfORaAUXXSL/NpprJnY8oQ2L8FHyg8r9DzXl7DW1AfQaObMDNSmUPL1E9Td7dfe
DYUuIlgM6rr8g6Ok7Vf8rJPP9kpHX4b7h1GGmYxyhvySZeqDOp3n2gpS1sKKE+mR
AKMSk+GauXqa1PsTe8i+KU4G+aiEHa5/QDVlOo1crYzS4dPFFLG0AnS75TFEpJM+
r4jN1qZ4joWBArUcSMuh8DT2XM1sD2eE308OiRv/ZhnzHlzeSkiLlJyl05Ynv/Uj
DWpmsv8kom3xS5iOtKnG65T6puK5zIT/xErF5Y3S0dJKDvZfqGUa8P+XC+GNkpGT
tSAy3hTU1MtvUsIxACttxCJ2KC3IO5Nx+ntLE/qAErijCPu8T6WQHGOViGXhyyNS
mThvdQNvfhGk4ZzDvIbfShY4C09acD3+ZLfxZwuoWBeFMzVoJPMGwlIHl0TcTgI4
3gXiNVeQMqiUH/JZxTac6c6ck84KXYDVexp2d8xW2LEGyFS+sjzQHSXtmsFOBUx3
1hckI9QWmRHOwb+AtJrizkCX4J6c9PUA21WuRj6LOrxzq8Y6FphiFU5mD4dyifkW
iq9uzOZchBMBySLleElxp/ZhxdMRFKF2oCELqLWA5OB1IgExLjrSnT7ehBUUB4xj
HqjcfsbZjPp3N8UPamNd+X2bBuroXmY6FqAHGl4zuyqwK5yLq8rndtvpCGiBe9/8
pZIX5cN0Bmy9igynT9CH87GMwiLtWUsOoFhUppKBo4lvKUD9O917WRZlB2rUcs9y
DwAy7+Op9zybbBSqfkfmQjxwWNvCWNGyOMo8kNwhDMiZXSjUQftCHl93smtROMzi
LY4LdJe/PZuoNR+2URxAmXb01oIehQJMcEQz3iPFn+afqPeANaqpkugqD0rWD05x
LA3Pgu6c22OpUOLYUCiyVcMyCUss/e1uX6HE+uz0WTtrX1ioMY0mUm3PbV+NzJw2
0mZBF7IWodxa98dJuo3apszUSzCyrk1dDiU05ocEIlmzsyRbc3SwNzH0MLGNnkH3
Iz7nOoaPzwjF3fvJw49q5OYE/CCKyGTyKkcio83SMvgIRzx5ZHaNDPlc0fVhLWl0
jqmvr1PFh+BPBDX5uuyaOc4obZC4B8I4D6VF7sZLPJOKzRaP2RmRWqHUG8lV1vNJ
V0gXjIVEnBGoOEth1/KjNZPLsC3CCMTBxOe0R3Mz5NiKyZfpUpPVQA8KkPkCNphE
H1V7BTh+/3vSewCBFt5ced0iMEi5bSA/nHYYZCZcP8rfeKSMnl/eMztZDX9XC/Y7
UAsN4U5BxitEFOwVCR/SCbBn8zGRQ8dbEkDss40VH8FZinJCovEmGVexGNg8MCC9
qmMm+YlRcYzUUcho1OLE+6dr1RZbza0IxAgAsAs8wNe3JjwcaZg6HpYWH7kuyk7h
3kzr/3ys15dhCZsBZPIXK52nMurHppYw7fQ97Rbth2aRqukp+oAucJhnJUUkgjfu
BM7L+NU8c2mW9dRrUoucFxxvhfCZvNznk8QB9o4Fcl/qT4Fht2tNdtRUh1VUeero
6bVJqoK0m1Rw1dj0O9jntnOVOdz2X927WmDGGD0zmS3fdOCw5vHmTSVxbYL34k44
jCH7lkIA0VLL05uIcvUxzlDbCxRFZ0TQaieikMnFv8FHb9ph7Vg+NKM0O/NC3kYt
EwcWWfxOIkcCY2/BDYhMgtrFUBqijnZNOBgziVx6IFj2F98STOzhcS047Dl17fgY
tSKr7o+5h826ZaFBYkVFI82B+vmXFguS/419l6TKRFNkSVOXJKFG0H9IzPt1VkJN
3Vb/XYv38G7sXMi886Vvknse1TZjxrsBiZrDFLhMgT581NplEJpGtqKn4cZDZK4T
d3LJyE0DaN0WmIIGfwCxUTia2Xz5EO81YxpPt/MrDrZeMzl61lVARcnlyTYKQNWt
rjaQ0SUn7EJMH9hdGZDyhAW2x7axS5V6b6gDmaoXj8+LbwS0EUa04LaFye96k8J4
08aPyCg3aJ8hsNTeQHWYPFHLCt/krhmHpg3+OIAM5gTUFjUWV3ikIsKt4A8cjh0K
+BRbGPpXL49xn7FeIjmXvgxk6OyUZQuI+6u4VqzbsuHbP2Sfi4oxg46f3wUopVsO
DMlJEGVjH7WmJL+mJDcM6mzYjxhMAQ2X9wlFddJ0tl6VpGBmo+7iiQY3Njb0d3Zk
QgADo90I79EPdL1ETX//cT0RVcEtel+vaCCrVpHITG9UfV+kCHu4PobAMP7dwhHr
SBADV4ASbrGEB6QvUwecFwc+xMzqS4tbyBmplGjPJXxWgyQFvEgQbw6V+le+epuO
DLrHlD48BOLNqwoibNSr/rQwSV7IU+eB0q/bDFQ/ssMfFxMENd+SielfPHDjzH69
LsTWFP8jvzV+5IPaAZlIunXULbB6YhrFx14egoy836rnEZ7OADJ/K6xOpMW8yJ5A
aUq1BnehYMiZD11HwEJRcJ9s1SYe9TItkXXlafA7SEC4yDG6KoYYmSlvjqSFMnEg
2jQDwRxnRvbQMjfa8H2JimCvoO7uoE02gIaI47DKMMSZ4dOFmmjQyR4fTECvBeyq
+ArRJBD38l2h60+E9RFbvwkD2TsT9fMFp2TuSE7pADO4buhX5ThhiV5UytUQxv2D
b9rbiQFwZwtcyi/zpv6dff/xqJr2jEbu3JX0ycI7l1WidKIPv0r+68cK+tMd0r43
55xrcptjZurvpx6Wb0K80jN+Ct08QE8ahqBSFYiLUdUNd7BZ5+DRjtNBJbe7rTAn
AgLsEulxj8ZiZxRMx50VezLqQZ1bHcLPOIqZUeo6RAxUcfTVMgDvt+dfE6Ux39l5
CmZqAEH4Zapx1ctDakagCtyXtaOmKm+XPW14/Ph/C0mbpkhSfz4sqwg5rv7/DQsN
SFGGGzqJy16+8deu/PJBd6urOoWYTIcdJo5e2a+h5BGXHskRpYKGRFvJAqJfRuAt
xe6rl4sIj/fJCgK+B9OevJjR7V3kzV8U1w8xA6+kZts85YkvSC1vDMKchGFe3mq+
4davboEFFrByYR2DMXmOKNlzgLFlEQThmnskrJfrj6kdXx9j7dDEiP+4CWJ7CCZA
51WKkAEyht1hbLUDVTWmcnubOwDleBQeS7TbG2jN1Ohg5CaBbaKRCBm7w3dJ4yVz
8fpWKkmYQArADhaa6RUKRlTkgjAtcjlMIt80TNzKfF06TQ9hrJp8Vi//CKJ5PR/+
obuL63mrLGOveAslQsMTIrPxs6RfACbjD2X0UMaTX2PCZPJ82xn9W+UXn6LJiV7D
Xend6biNKPiIpKIX69mg5x/4PEYlT+LAF9UtMTF5WPEN3rtQxjjp+OlGt/3XDCnL
P7VpGLhJuK1MtlyHV4FxPqYx9ENtGbWRX9WnRdY2oj9m24ZeLiz/hBS2lOD7/mDS
tZXN6wLvh77R+wfu+WadN3rrAkZutKqW0PnkzoYvFO+/xX/6REes7D4T5pu/rtOe
7ARku2Uz54Y9BgZij9N8cuzt36+gV0PHN1Sj4ZKVnmcA5m0jJuwZGdIwxE7suWec
q7WkXInMTl3QEdIBDmMrre6lnJz1f61rdYGwiy2yVUOTvPP/R0+msb6xsxFiUKxs
Jj2EZJIGpJmpCCvMN6pH4seZf2no2lPz7FPwPFOcGlt4oogNuBHKync7CLczg+dC
uyTts7p8QAuT2SKIiPLiMZNXvc4waaPuBD4FJad3cxclEoIF6Bsjb07CKfzE3507
wPehXZ1nL8V/QJl2PXXoknASAmT+fyrRM+5d9BmA1QXayEpq+9eOnTBFPg8YbbH2
d2wHzuEQyHZH32qznCM/A/RRlaGhcsOPqBluGSOuHiw08N943QPnEdMpnWL6zGrA
cI6s+3DTFUF11hI5PfBuL/cjMz9Aea/BaxDlf4QeCpgSCA6CHRUmBwEv944uMO7s
IY7BewO6IKn2X4WbMTIQCc9T4quFwHA6kfVPlEt+dlWH6l1gBx9u/eLPb012i3EW
x+fIpM/xW1Vlh52mMcXEsRTEeMqW6E0gC4sLaRVvLbh1vnPWqyS9iXUHjrFXoSdH
dcKaAFSdqzPJbuGAk7s4sL0xK36ofULsCdd87nVplpqR8ccTgwwqj0kjjw3hE/ax
3EnIHYCpBZFxMLH81sKqhpFHQ9aP7eSN24xoLWlFGl0zHBD0n/TUqbTamzBu5MPF
SyopeOBpn4hfbwFCi8Ukn7E4oumznj77YolPU/6AVM/wnLyu++tUjgzhFAhjV52w
q8ZdO28CwkZirIod/ciX7avdkuuS8ADI2S08uDCp7ywzGSlR/xcjDUM4B1vypCQp
4VNc15UEWChlc9AngfuS1j+2HT4zNtBa/tl9bGfbkw5Mr20BOjTjmiSPLCUttbsQ
5orjWlhaUDsgCp1mcEd5hDzq76GyVkTn8g6bwUuaTHm9uQeXfjfolP+kscR6gLXD
48mAMd1iC7D1DxNOB7la8+5pHLlwq9OjsH11PRrG+dRbvupyc07VZZkbC3lgs4ic
F5NOVosrdtzSbnzfyZ4ANFIVXb0ccuR2WidwLl8EDvYj9FTn/kHFO5p9kSRBGUMg
ks4TmvEPBove5otSlC9uw6zm19Yvh133vztkTzTg20OsF95Z+Ul+QAZfCHNLJv9a
1NzxS3oLge9Em5oE/Bu5m2bLq7HUOpl060f6PiHT328xNfOfmy/frQwqtjpmafTL
0ia/cLHn/7cK35D+o+hFyBVj1XrOObhi3zk8nEVYLLDk7v0x+9XkdsHXdzHfoAj9
6rdPRMU6jiAkQBZBXAXDNM7xFJd8juHE5MBTDvzGN/6Ktxj/J1UE1b28UIUrFuTG
AcxiIyneHNTYGkLBjGXACIHOfJ+bmfcC6CjOdKfho9jnGAPXmFS7XbrGrOSdvuLk
I0924v4tkaule5OyRhTdPfTKpXY+Ee6pYrkYENOxofSvsSdxIJ7tAOBwp+4oGcI3
Kf21guIY4Xfb5hkgl+TD35vSUnacRZjxyFFIgZCIDaWVcB8/llZFPipt5WLfIX6N
Jq8PB5Ew9oZYkKhNCsEjFTangkTPs0WIjR45A1ryY6hrBWBCWWdaYoBxVxDBARdG
7h3BJRsGd70Q0e0FWeyiIisiXmE/xr2EknH0wVmjtzroZ/gArDnMCco+khEtOMb0
Wmsc6YjYvDlph6fkc9HpIFq/JlCTvmpruTzzIHrHzApACKqcDp80RtCH4xGEI/uN
ZFHeB1J2gqyMq9LohWeAy5QFTMaLfgGzevsdxUKric/LscoeO1geoX3VdVCIeJM6
pp6840nD/utEwrmoq/PfcrJ8Q5rktbe6jP/xRrMEzhVDJSxffQkUDIGD18b+SpwR
B58is+j0ykPB7F+/QOhdhYsgD6bo203uNJsCqWrxKYpnKYzhbtFNoSISE1oiIooy
aAVyLe/UVTugSxcVaBTW7TInVW3iXLmwJM8YBRgOn8yAe3gaW18fIg0MStHv/h25
9vYHKU5LugT2GuBBQGa8T+c6/cnyzKIryR8NrAiCiUmdXz66uiiTVQN+5c/Hjdlg
St/+UTNoH7lBSfzUzdGc0mIXHMFwjG4z4Z1aLrHupva1aLnTbvTbMPE7rYfAjoJt
xSbkRrODzW7j7wtQVlLbHXesh1ZTqPvWWG0+6Sn4xw60IjSs5rounHor+unATq5w
II1gHjqvFuCVBALHiIXf8WDtZiO2YI6sSjzV49vm9xuEuqrcc8X/PNZX20kDta1f
Nkave86txmmo9D5WcuyIaUpVV0mhyljwuiqXLU5sCA1q65CUbo8y3ycG08jKtU4W
Kgg0Wx0bg3BfPEEehHlxB35vHVHaSB4EtBtayTt73mNUH7ERxhjMKIDzQ7IF1l2R
M84R+JDQp912vxReWEayOY6dURaEKnVlMpz8mBxkoKOurKpKFbrV/i+9PuK5bKN0
eeij4cKjNhR2ty+syZWBQN7yByEY7gkA13UzLRqofZj3HLpv9wvFk35pgM8hfYKP
BuFL7qSKzMhgPMJJwY7diZJL72WRdCtQHgmCTZZJADtxL3dbjTOhZAT0sAJVmuu2
pXZmTHnstwozxuH6Y5mEm+hQeuvMRBmyeoblLE0JwVuYfcI6PWoYxfFR4K3Tp0pv
mug//EdhOGndBSw2JzBvqfUIfdR5B1yr1HOtHPdEECZfWexzk1+BSc4qi16bNIY/
UNPchfYj5XdOlKBYJKtq6rq8Cxb6dvhUfEm1WsAeqKM2NpQv2tP8rtV7X1m3KMCe
/rd+WNz+s+vCC5T1W2uprXs84fyhXkwagcFFvH9fkzZO86Za7U0NoyP7/by77QMK
0eKgcN4yJew16gurVkCA24yLzgv4FeJ0aS5foyFrr2grcQWhWPVv2i7rqRLGYrXb
4KhhA6ksqTjcYN0GslKKR0eGZhipsqbXsAYKl7ZhI0DTPUnbHRa73xNX7ZrYI4Kb
zuSufRgw8sm5acqSh1IBR63wg8if3TvdPIpqdAjkEtc=
--pragma protect end_data_block
--pragma protect digest_block
w1SD5HFxUPsBkJqaqk0Qi63dJV8=
--pragma protect end_digest_block
--pragma protect end_protected
