// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
pbKDFXKmR59nmcljRcg0sjD4tWwHEyx5YfkaW8KpAU/5nkPU+SgTf5+VmheaVZ+oKrTouvx+ZS0z
PmY/30HiuPmbQegu2mIgTAcpByaHfrUX3Yt+Z8ZqAdN40Kk+FnEKb9OakqPx/xN4e08RgHaT/PqU
CuISW2bn4GbFK18qqLBDv9bsoZA1Iw7kRi33cXUI+2vqKWyERU+o8pPag7UObmaGpRWJ0EfW1Ne2
JhIftNdWxt9CVqv6a5MbMC6XKHM0XTH8mAAuy5o088vT1Jl+ITA0feUGz681bpPSuHkP0Y72h0DW
7jYLJexQCa/yjv4zygCND2YKmPk4pgvNLXqMXg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 13536)
2druUl0ThDIvWmZx0zgBkNrsJ+frtxVFQHBa+7LW2BLpR8GOlNjXBzF8HDVeiDJl0EQFosq7PKFW
K2IpCYAp6y0yd04K+ejEjvO6O+tBggTVRURlUjeayJjXEPttRQz60b4Y2G9/AovGguYLHDyw6vKc
aS10ILWvKtBWQ3+wS/tNson00qWW1w5tlAa2PrO2rUd76PBozDlVI+w9EJyAauVzu6bunvSkerYn
u6jxoci0uBtK/r53eDhp2joESvwxxmiBupBSYyJhLdwUCcvMvjtH64Q0Yaf4xaxTuCDazix38lE9
J1yL2S1RPyzuX+NNN5LEyARyx4J0hHyEdcGAIf+WG8s+qkbgIKce4ehEk9nJzoZppqRFzN4XHlg1
96baipb78MsEf4jrUUMOH8eX7ileexdsNu/W5H/9ThzzWfd6R4+TWKXsZph5cGWoTHCPUfqQ9W8n
ixZjtTwu9w30+lkqrsRyH3TIcCvsu7H3mKl1rHn1quJZWPgx/uH0UMGqUdYA6t6LsXUbbFHywB5/
GBa1X+aEFQBxNEMH2NxW2V1VRq+6hc+E62vk/HZNbWDomxM/R58iROANkRwI/ChsKhTITMNh+LMM
LBFnL3sEgKqGoV/+s0aqhq8c2EQhtS1IJSZA8yYnUPOfA749NkLrAVmP4yase6p0/niqrzGT7hxF
jpEKy8v6iFydeDxhZJ4yTFCrPpGn0t6zWEA32Ehh4DxixUgbUjJzGYZEVsBP/nkN31waLnrrmdt1
MARr40a1eL2LC0zwTFQtchZSbMcZQfz27ZlcYwoLweHL7FzMzrS8J/6KOtl7luiDaCW4exZYlOSU
rJSdnWCodGKbKgAiu7738cuMZTAXHCu/WV3saJQ/rP30XfAUhtlBGhg5jsm5YGo0JCAeVCfYK+YD
owZzuUKUzpXqPnXyuH6G1TfG6K6sJ2wAqaVwWKgq0RHa3xtU3iAVSqXBmixWKvcZvO4wLcxY3zaP
LzFkmKVSyVPoYxhu7CpAKXr7VPptmn4u3nRdFiiGRHustV/vlo5tZEdv+XtAAneCAn8A7Gjnh/ZB
ryXdw1QpnHy9zF2Wbw6iMPnZclcuVhJM37hbDM9Mj6Ui0x7TU6I9TQUAjQgpa/5p/IhpZ6QSsPed
Dqvp0UjiWb67S/TorMjKm2UZziKJ/ZxwFGjERUho0OpZ340XjqhK5eYJBqRF8Zsx14oRJ68Tqyh+
ikYVQZqc1JXgmg57bp3nt1xiUsDnIr2fW9g2ayui6lXpGc92bifdTAysUlrVHrXvOvT4uQKvKcdl
1vsXDN0mK4y2IODFsKQp0gvEptVfw4NPplLVRveX74E50kmq4eR/zVrFGc9WEnlqqlrgb4dwck4A
PHt8GgxXbZdPvqnP9yvFVQ0cVkh4my/Ss7EyQBCkpq4qxzNVAdi7DmRxeE/0I1f69U/SKp0mcDYU
Nr8gNyYyF6wat6nQl+vIGAw6oVT7eum1prYhBumm5EbukjqUiPQy5vMf7505Xkybsq1fN6n2w7JL
aciRd7ifePpKoiLXHe15fBuRenLAEGeK0aniE0jgTyAZxy5whJ4dVU9PthcUDlMKjj9TrOmMrFFx
Fp88nzlwdIg912CthHzhri75P1xSxSvMarI9qbNJtHJOjJLRe46/AgybkPyCX7P0yBQ1uf/TuIr3
y/dddLTqbjkJQi00vHiNUEgVbfCrPaEqrFaEOLjv0TfN4N9nTGdNTeFmj4zxRTyebgTfle7P9quQ
htDNEwk5asoDHBGy55BeX39uavHVqpEzaInQmNakQedTXb8V62913x7c0CcuO/4EtX2du4HosNE3
BK3pUVuVKOrdao7w4DH/3/sxYyKsGT4kIWMha7yn+PjXGMyM8GvlkXqArRfO/PHfLvhyy1hTrrov
8MCGAqWdgaHQfxfx/gZrvhIFeDgEq7oFc6YZd76+bVZuT5px7KA9uO3+P43DZEGJ5pkijHrKdilK
wWadMQt5J0Rg3+1U8pd5Pq94jP1E5DT3ozg3DMqcFhq3FfGxsNjHMWgnmGzhl0Yb76RuxuZP/dd8
Gnu9LSJr0kvI6TzGfLTBj0aOqK/ENuT5ZeC/s8eL2YVoHQwZ7zoAyryaiMsE4ywwVFHIITNpsVPs
d9tlboi01IBQjnBjUVuE1e4a50QmgYpvdYLnQOaUzOZrg1i5GK1OJRu4qB8cvuwAMx8jJsi84H5g
8ZgM95tp7i+JZpG4W6REiW8LSObetvJHsidUv9eQieVRYvFEuRJhqsZ1Wfx/LhH2LTQypW4ZEwgs
Lrrlm0ryjBhWG74u2jZ0g0MC968wjGWVPj+VHf9pa09sM5KmzzVu7vL4JJReO0fvmZtNAf01lGUB
D3YymYrPXmYcIDfa+KR68e6bLhB5KyNIJIadmUZkEXKvJjIgt5z3kcz+7VZeNIIfgkNorsvQgWR9
bf9wuNosJxM2K37Ndky84UIYjVgWBD9Uptg9SOqLV8nNN2RxGwT3xV7iyKN2ji87BT+FWsr3hq1F
jEFUhT2y4UiRzh21juYBZVryfTyJCOwOPQT2U5EIyNeOTlUzBRKvfzeYcuS/L435Ck+LHZKaJMSt
cTT7pI+/YRzhfzcNKkCrYHp4prwikINZtWz1Z/bv79aXwd6SGaFT8dijjXpofl8hpch44M+R/Lfl
lXP+vh/rV597i8MYUQ1GCCMzyOFJkYDS6ip9z8NbPR5FnXFMS33OqwcohOVyfVVnuAU1Pin3615E
q3pE1I0J6tquPN15ibLekWaDHmNjT5HJaETWRK/fQLJsZVP2mCHX/BAcj4khK23t9YLw8VxQna1K
2BO8t6BFt0MblcMVa7x4xPsjU7FR4Zrqz9VOOCjyPgymg1uEsVAe45C098883YnsyXHLoaxFn+AP
7kg8F82xHWWbmCfGZnZUljUdBQbX3VwXRoo33npY/SxRZuWndSwuuowX5vN5vhSrXWUrnJr9eHGt
60SdPY5/PfZaUFUQ7r6JTtEdVhzyh5NAaTdomIyaDEJuWYybwlVErM1KP0Vo6eYz1MKDU8YA4Gpo
gpQ6aL7++GnCZ+uaIt8UwnTBmGiXJo6KyJGpTDiMwmmch4D1ydsEN1rCEBGfv3oglxrvmVUsWXRa
pV4j4tkIMybKr62U4tAcmS1Oq06OJASSQEzAavgNCZullan/OtlxnwfQIMKeu3l/A8c0BOb+kaa6
HS18FyGpeb20apjY1F1jKJWl4Fzb4u8zT13UsD7+jK0ap8HmwByBiApe4ImmsEQECo7WyIq+x6nu
PvcAZra8YSEQnWGDuzUGU8xU0g2K0p6wv63ZHcdwcjfI2bPZJi/m1Pr+CrNUSumTwKwLilTvSjQe
ABs5rwMeVPsG93jN7P4K2tW7t8gx4KqnLPjTPdRsh3hMa5zHDR+pTVENDE+xHMv7HYWKvGJaQGGo
z0PGU9zl2YXnlVKvS2t4VGfwXG6jjOLPLi9IAI9Pd1W3p7RULjgYd/WVNKKFB7LwNKA0rUKDrBz5
nzqKEgQ1RsviPtpkN+3VTZqHMGT3uNzwEKewmvD0DCLM5Xb+Hk5nw8WLjWNM59gpdA1FPRPjwC/j
TmYQtpTausIhYx9cwYn1DY++IdQ9NAYz6USq/CCOCahx81V2E+zwyiBl9oWZxZvJ5LCiEuFKHIhH
sqC7J1IGmCvA5/9Ao8vBcSptKEpBPcY+A/YwKC8YcPUrF8RPNBCyNnx0E52lyy11haMUUICCOch4
KfY+OjRyzK3l+T9haj0UOcfdjUSPEsXMYm2lvyNJkoER41ms9wItsWr0e0VGANTq6bCLUhI0Ra7d
mcPZdrdIm4QvNfzNEnRXLuFmX+6NlJEc+6MRE9F4XtAd46RaZcUP/oBHIzNxNTv11ZFZo3n/UI1s
z5cD2sVtg+b2mXKubYDk+CHEelsapoAJWYNy1wf2k18vIdKONj2RBIt7++iP8v4GWMmYnUs+ZSly
TO8oIhZyr9AXbzOJOM8MHWVC9IrTxg1JXcGmyccDbxJBNacEUdFGyC6AyhWGva2EzPEBWL7vtpJm
sDWMeb+30DKm4DzhPXN4iXpSBKgQWJTL/9snOFqtMR9IgfX+sHUnYTnIl9TshWCmcvQL0VDfMKKt
0Chnhb/GVhEmNBSPyFg4c8DxSUiwUuH5UP7pBl+BHpGTVtRhFRFj8uYHQV+G9WqErAhpIf81eHXC
Tz8jsBb1myBDb8Uvodd7y5+1IJByRN4lWGgQHYgv5JC7+zaOKkJyuMdEi9MlHKCS93eZA1X4XMpf
cn+eJFDi48H/03q5Ss5eTFTRGMCvg/uwbDgzCO3VK4Rb6FQ0jaryOJ/KrYw4pxdzIEaD0jg9453d
vbGU/ruTsYyn/D5yavJkxQet9XMn4p4wTPlQWtrRy09qsIzSI+98sOlaeVPeJxKKmhokx3qxwPzO
fbhhnv2q2Aw3bjKM1JQ2PncbRJVGb/6xtq4dBXO7/2pmqlHorI/JiJ4tSTV6dBJ721iLw52SGKKe
mw+SRZabarfbNLVJgyr1lf8xIFNXOcboiK0tczuQpn71dAk1T1saT2CS6QrJsknhsE6JnQ9LgwTd
TB90+WQaILG+whSScf02ZaAKy6HVC3KWssGGVt1TotJOipAinlW/7bVcevq4LMiWuXViLWv05AoA
aXljXG2nE3MPd7lx0zAFRJrJjKfgOnnGTDEzP9wfmHzMhBEOcPNfEhd3Gn1m2nSIHh+PLNVPsmk7
oJAkrzALaTroTajE6RlKUjJJlcDVy372CkIUueSzJwiGEV+LZ9MCKQvy12j0w+tyZAlWgdggKckA
9O9DLrNnBeEx3FT8JOVZ0owS4VR61fJ2g45Cn2N2oJYKN5SNyAoQEhtTJVFCPnzO1ymkP9GJj+jC
hkU7tZYO+HBoQEASJDpw1U/3qrWC7Y0N7k4BCFOrZF/vYHrXbtfM89WzLI6/WA2F3NUSQXzHOTOg
udoxtq0TF4cwjC+3sAXzweGhBodzmu99crqzAeT+hZS2tpKQXJgV2v9F6JotFC/W0G9KJcEB0RVl
Cl92nswdXiBTAAS9l0cJ3oEL2SNKWdxGm8/jQTSwM4frga1Wg6qw5o+foFTGsXKwE6xWoAih+QWC
zKoIM3r3I+y7x3etdAm7tuyKYfNWeD+XUhMasD2t8WD+zDIbSuBfp1wvQPqe+ClsljxJFuoiXlCF
Ur70MCk7gorqbLxMcaka9Ancy7wDngTleTYFkqsGIF+hWlhufajgjU80WoJtaJYNdg00y03Cc4l/
ESDTzGFjTeHBNZERy8NpyG/FzQ+3+8BRWiInjw2Hw0mw4GqjE2cY7d8jyKnbHVKjwM20NFq9v9XH
HosPZsbVPS4BUs8bYkPcuS5FJ/UNrLjh3cWHu954A6vdkTL+FHQG6HHQ4lmnuHBImNh9IUU/AG/z
ECgr2q1wg2uEu/DtzkagxhullO3u1OQjK73Gt4BnsiTWeRUUYkcheR3EKa5SY/++XEC4LIvLgEwc
zuJElQ2zm3hQB4hV3oZRG7dT9+JDyBgs3EFOisq14HR4iCPHzZlCMnT8rjLNW8nukTZM6VumGzRE
mn5YPIQ0QCoMlEeBaQSIHiztXjVnpNfR7jzXMrPiFwBMFAHgAfKAntOvVo1J/4g/PUvPLAmdtV21
kpDAlj3GtwjIm6gyBa/EcClzXQUX42pz2V9C09mN/9YgSdNuaqp1rDghiZRiix4ccdMM2TX5OZ4U
4BtAbrcFXaphuCBwjCb6xXnQ9cbpUrhpOWIcD0TbFXDcqJZY5W42IBh7E01bmdv8ZaB5BNpHtwnH
X1u+1nq0de18GUE/VEp6lofi2tSipBPONqtNCm3J9pO4i1/Ab5SUmElfe9XfddyYGWS5Ikg3duzI
tyEJYsoOpQ6IjBMP4bidxOCA14z87oXKb+l2y/FIBvWImVY5t+47YpyRur+M73rFULkIDTgJQCz3
OOpa/5LMlujQgAyE9eKeHpQ8I7/141+LTXHIk9tjDD4Iw/VtvsIR25Om28/RvVDiPfolTIa4hapB
No8a0+VNU6iQfZ1nxYFWdokKG3XMuNwDfgj1Z3yzh7IWk34l5kYY8yLUi8gK44TJBabPuVIoB88+
pliMp/rjYrYVazaruSvJTXTFYCrBZ+wnsdxZD2FJ3UgTG1nBvRRL1qpgJrODDZ+6TssJM3QRZq3m
On85tOBsZ6Ptbjyo7ZW4Qt7JEB+rXvGS4Pmv6n3uoUIpBOFrcqocvVAO7TwrsH0m8zcMJuzilThT
9ma5xF8HvMQSWkGrgTtu2JUumczMl387WI3y1ojNAKAZOIZQqJE5LL2ej2VR3qJxM7mPzyo+polt
qGmAR7QX/u6JS6XMX5fSZAh7VgOjIbAfsAz5WNZQPdD5vMkwtV5pGcoPCOFU08D+1Pkos0CFdl1B
TPK4OqJcLAbplU8WgHWm6q9ZIs5dxnlUsvtu+1q3kzuHLoQF/8AjEpg/lJg+XJtjHi2lUDY7x1Gd
xKXkmjxtcLMcJNnzXWRM3oXZC4AQ/3db95NrbOVcw+7Rrvyr5ojQwMyCs1prmsyip1ZjlB3dYJIg
POZltLYWkGszgIfftWrV0gXWrqT+oEKpZDSTgS36PHukYKuorBjrv9v17CMdtnhWTkktPcKSFFAU
eURQ0C3ueTYENbIWDUIl4xohwr7onm2y3TVBWGWBzgQp6TxPnLfFlBBHBRt75ohjNnssWWLgPAoE
t/XQSbxAayqXjmKHu9o5P6BEK4fJHQ4pOzu+JWGqUFRVH4vh00rdhOleseynebU0Fcn5fymu1ALg
w55/chFmL/7YY1PyLzUxvTD6YfMw7gnAr9tbOmrorgBRJke7UUjJ6ZbaRY4JnOORSUZC5jztfeqy
mL4rdRnSVUN1x/zH/lVW7+UFRzimqMa7sL6vYQ4BVbJ4tdoo8d4L5FqwY6nCDz/axzXSDbnVK15+
tsZf0EcsWqb7n8uNOVCTkNgEVS7siQUQ8bNyT6VICQOXXK/s/9NwobY2Q1076VbmEdubwgzosnRm
7JRTHjIyafD0N1KN+5cNfSIooJpFboeOHBoJT2Gx15CLjiW/uZ6tG8GQFAbck+AuiiPJF3dEeeMs
QoRJMGMlhtSeUCHlfE1VMNdxyWjGmB6rDcvHYpM+YzIqLzn9HKz3IiNl6trpzXZgzAWkx3J75XmN
Tsr0NJHlaCFPu/pA3Z/UcRQxbAVOEEDwJReFkBXElUv9zWdwVL6aMckrTwoRb935CB2iAFrSoe42
FgC+ZRLFwToEDxzD5rwuX8+UYCluHOGwsF3+EqsSJYaKNUamaj2uX9WtBP3ZmxsCIdpgnPGhTcBc
oYi3GvHX/WqTFt4qCUBB3XGacn7JDFqRTzLjNtYAUNYWlZVGv4sOq+ZVw0n8Q2uoeS0CYw+RNWID
TQjzqX9/PZgoj/qDwUqWvOsopmhWJwOs07spxG6SCXKmdsKNgSoDgyhrQ4QFnYFHQEfuFtOiU3ld
GnHdL8SOPnocPdWTmzO/sdSTTLkK/ji2HjYUko355hCDxxvZjEDW4yKXLFaK/5raI3jJR1JJJnnQ
/ecgafda3zOMBdKfyadobSD++g32maCMdL/d+LpkxCOkrZkyH228RcPxYzh4Oev/rDGoZprzXK12
D5i2kvvyExx44hDWCT62WQG0K8hg0XmhBneW7r76+EBRF2Cp2OTuH+MxdjksAyAO3uZ6szK1gYFZ
zjZobEdxsaCmgFScLhvCJToGP/T1sLmBI6iBOhVLQQVLNeJc5R7MjPbBCCfAVTlasF7A9Uo7RbiE
xCCuSbKnZHkP+bE0V77NkjvrnBdJiVMA89SOYO9vGgSuVsFSiMQQ9Y1lyDGcbhotfRbt9YkY33HI
v2dhSBAN0rqpPkrl1SgOSnoI1v0bwx5y4e4tI/31R2gFAcDmVvc6mHITYwPGeZM3RcxjL9zWei3Y
zQSYXXVsC/BWajnSbP0zTNtFDbRcsXxTiKdX5xe6cH2o4xKMfYRQt1H0UTtRVZDjeDnf+Qy5Th+Q
e3aWs+KiHiigXSvPyGYbxvIgY8R8UT8QJx36n/WsOolSg3aTWdMsyDFehBTDbgndNskHNenIcT45
0uanFqyVU67V+vFMuz2WZCRhmgVDUccmS133ryrK4R/ilgbntcBPI7pBaCu/ao6h4L4jBIK7PjnY
VUABWN5X4tnpH7FO6ZRCgPBtsHDb3d7KCIguUYbOFNecWqi2OeuaiozDvvjAGbSW2yJIfnTxWdZ5
/berfxy6oiwXndX0h3Xtnm5FCrjHhnCqAiZ2h6MCrLZUyjIKgaOHEa4tCOO8+nUvMoAET6KgeXoo
+dQO/GEQ0v4ovcZTBO8kQ66Gib0gcWW8OH+f4bQpiRcjw2RGZgkHDyEjVY96smmWYAUHi0rfslaC
5dzmppRchBfWmiukrjaF2elsrIcy4l3sbRTdnmrtdqyTMaaj3zyREXv5GS0O1MnlYnIf0z0ALfwD
s9dESXQuGtaItrzLTJ3pnMWWu7WL2q7sid5rc+L471ZTe/6R/mbJpciCMUt0WmoNDoFptwZo3l0O
FbJ+24u1FtNOIXnxhfp8lZ1SwMP5eRYXWW0ARYjF0dQF5FTJG6sXb7atY8p8f9i9a3HNad3IZxpc
vECtpxldb3+0nAx9cM3k2IYbKk6t/+7IRchnPWNu+1bhICiQFerc3TnNeEZaWpWpx4HD6Y2QPGn8
35THRGpVm0kOY001TiQ4USTygphH+gl/A7eBjyoLBiFP4ttup7RgwG90HxSt0q3UPm+5xDG5OwuQ
jb5opSGsv5/eGVQ5oyYkk671sWjH5whoHHRiToewG944YYgjnqTw5Bhq2Q1t4lx7Jdd794c43CWr
QdFHeF0DZXn90A54j1M4oYV+Q4RQhul5M8wIgRwf9t61fnlga7KXm5Eq7lP/k7g2w7/cGcsAanz3
Wc/T77thvLjiGfMKyCO9sNnNUzr8kxMjBMDAYaZWHgO2l7/wftpjzW1D1ggz1Mg+ooSQjeVu35QE
jdazQso67RROfaZHxfA176f5sASG6lS8zdfGn5RYbPySu2Ngp+SSD7qhIKuQSXipR+JkmraLGhN9
EfdHdbLKTw4ojQX82MVOK/osNeeiH5RH6AB6sD10HKcuQCEQfP/BGC85lFoL5SZ5y8Fh47jafWBv
647Phl7R73d73XeBaqrnFS3/7w4Vywc+NMQCHxfANsQ/Hn2nTRZXZjVy4rXBBuEvblxnYkS0KYaX
l5pF2slwtbWys/wRLl1ykaz3lpKIaVERi7nc1WDu9UModJLN6Hs2XvIQOaEDp7djAqxb/5900yxY
d35mFQTll4TgYoi47pov992wLrhsc+DdSR9VOIYOjtCtxEqNGYNA/+y6qVMkNcwmqGqx5AoU8nSd
C3OcYfXAfxIHDtGMdNmOpnar/HytP8qqWbz4RF43JsfrCmGgmijJz4m88XeK1o5V1F4M7m01yTOY
MmS745au6D+XXnP0wA/jKTKJWxJJpBjv8jcXc+Rc1gP+YQ17UmlogOstXDQqgJYDVWIuZLNAdT1N
b3t5aJevkqR1yyiYm1QZNQuP6V4usGSL+8JTVIVktbeWKJDs26ZRjBkJ/63bUIRc9nA5GvIy4zWL
ZcNedZvEKg9cyl6M5qMJ+jDQDQfDETPWeCrAw9Q62pNiABqSfSGw31DU91cR1OjjwoCKNXzY9T4x
IwcHdkmpRBPL2w2ihdE+b9JADcVCkvXHik+g2WmryDmMMImTtGaVPAz3u9bsY7CaesBnvzlfT3Gd
6POk/dpaE/1VzCfcfZRh20bOAmBFbTEKpKf2st6MOX34+GYbqdRMxgNExeTbKUJVVxxYrCBJFOX4
LoqOxbnZM8i0WbkLKOT88OHlwM+qSkYy09AB+IznNspAYuhP/FfTNJ6lpIJeU6Zv4ZDIdxJEFi1L
VllLickSI8/N+/JB72pvG/mCHyIr3H0n7/lVWC4VsSYsh0rfwh6JvzGuI+x01t+TU1qwb4DfeBOO
9/1onYsBqNekM5WFCb0w5nwrz8mAD3qi5xYuHdNRoByoVNdXxEbQcl1vJOtLtMyOKffIjLbtDsC9
v+jn3Art3QnbI2sUdHu7e0RBmBjspKcEH9zp/NwGveBfMkJJqnUgO6A6o9AKA0GKcNSI9CakBJfN
l0elDw5h1LR3E1kvshppC53uLQifvykA4nmM2wo170Qxz2NI3X6mwFFHSznvmSkCWVxtYsnb6uKk
rBFop0LSoKErmOMdxRINf9C1vgh43CpPA9P0j8DLHSlNaYI0VLPGKNMdoL3f9IaqRLY6OSpiXENX
8MGq+u9s7+doaBrWVL4mG/6N/cdzpKMbTx7A1l9wzSwzcK271WxlAOCmIY45x+ChpNmCE2N34Chs
hAC3+bD3T3EBKPdS4+gvk3TOBGkga5/tuEEofKEk+LnI7XW+RJczAwE6wA4auTLPd070U7D+8qUK
4/x66YV8rcktrPh2lB1COqMzVZmAl42zEwAfx+L/J+ldWJRKrd6zwipn2sveC6BmdIJIXKFfchn3
gtyJMjLB8cuTLfL/EumS12A/T2QGW+623TxHIAHn+3poTXF+9XGycozTpGqdM+RbjqUpxamy+rtT
0R35EQCyGFIwR6bkBa+w9ZUrwbzDKUvVcBz2OaH00SKP+aVLnDuNmmCVXzaY3utBR07oxwMPoI0j
89u2KXbzgomN6v5CmPos+LVSWFRiuev3DI0W96afWVX4c4/DFXAeFUv5KrkIFK/s7SYax5wHPwd6
eSUzOdgczl2+o3DzqoY5BB2QFYxRu3o+7CnciZFNH4QXmN5OfgNahNA69hjW01ildxR1QMdW8qfp
UQJ/JYL68iPrF6nCeOyWxXy9LhxkfBQivEVS37H7/JDPJ18r4uYRjzsgNOpGBhS3CHERdiOeRUyS
yApKhe0GTuzguldNsEoO2EBpwpSyTH+7Fhv44plBC3c0yi1SehYjnVWzOltFWiMFeuacPtJkkjtY
xjjRW746tVilMJ4sgeAjBjhbQnI9bGpF7jW30VYWayUhX0i87R8B4U631VNY/YV/U6zwoKqQQj1G
SwP7RkQWKcOmKjrty75o4SDA9jJHm5+U62aylNNDydFzX+VdXoeYknnlmfM8jHc1IfjJar3phEUM
k/CV96p2CffRg1tnc5KJw0urHj9X1lEcedblIANa5C+pBn5y71yu3tFlNhdN/uoKgCxRRHhiF7kx
ZwUoOiFhjxDOMmiBrRDc5fiQPJs/NC0nj8eFvVCZ4P9FQCNKkLmv9nmYavMEJdzZU//u540q5I08
pNeUSnhgW9Ex/D8Iz14WjjbgenGzPtt5aLcS2BWRb2rYl/MJpS7D4ilRnq2zeFAPoZ1s87JiAYvW
70PMK1EnBMqmOfV38VY5eVZn3j1ezBQDqVXETRDfK3SfXjAvdl3x7SGywU2YBigUDLqXssH2QHqA
rn+CpnobWEsCzyaqSCHIK4mXgcmkZP6H4WuXQK7+AXpCZ+rNEyaQxz7GH/Xxl1UC8A6vAVrkYDsG
affDiYgIg6vbleXV00Cy3T4By1pvJvdSkaaZo4Qgzh+JiSY5/d7dkuu53FPi4Y0p0bjpVB+H1JM3
jM6sK9DveC5Kl9tyabjHfFBKlJtoAYmP7ROyZ4Dky05/GTYsr6qRhEf+uuwemsOVM+NUmMy5k/nM
nxepLHaHvRwY3fGRpUMHmHnqAJi0DzIv0OyyGHKTDguHMG1pj6RHBcf1sgSgU8HDIDqKpM/DixBX
yImJpiWVtliznSfauiN0YCX0GH9oVsTkH48T5BJY+wrnctB0qOcw5MF40pjf4+12z8YKEgpUToH8
b5e978XpifYUAHXNGB0HybhtgpuD/p0CYUhuZo0ycjDSKOGAVBQx7lJF+dtzmQ/h404FigvXubv4
iZx97VFd2PQ/KhYpgKKnhbTTkHD8ry++KO5pV2k32vGeq2m4DNBUJvQVphez0Kaw9jZ3LFEDEyFT
TswpStQWX5q7HIlsPB2bva88GhhLsz9FaH2R2aSX+AnG7xkYkOASILeZ4pmgniua8pyF9n3oqojn
3ZJgmKHS1cKFPY9XkalHw24RJYHxMbIrRYVmRrg3dYQCEEmr4vWeQc4uclAhbZr8gCOzvrWUHvr4
Qy4pzJE99yafh1vlrLgtVw+uDBB6qo5SsZl4MQqyVG9ACtT19WpcaijUkj6qwew3ZDOOAPMLGe8S
YKTjcA4HXDwxdwmTInIm8K9/iDEkHcCfEgzGjTF54LwcintadspHCWNN6UzUxSvZZz739/Z6W/Hy
AeDqI5WjAOPL0FyMrO6Xr0z46Q9v/+M+aRevBTPsiSC1XjXFbABT1aEg49/380OUytlTGnkDpoxN
wqQS8uDVwDST51Ahy0PtOX7lgEzr6VdvW2jzFJbK2mqoPTguNTYyelukwHLYi/AWSRe9sA0g78RA
EsFb6Jsjl6/hjT09UtugkX4PYGsf5xVnaBgSULagWlesZ6f5VOnLaeGj4QRm4oTu2UHUj2NCwhV7
dGbjevRzAK39zlzmFAHHcy0npOpDEhtSobG8UVab+6JuMP8g0E5bK2VQ/Ao1i1ePWQxIDcAxCbw+
+LvMJ/g+Zgq+t7Rf5Yv3wM/sLRuFTjLJaXjMzoKMYftdhhIShwcI+erTL2pUy21Am6OzVcdNDB4/
B6nOKikGzyZrig2MnbYAW6hiQGsBthDwSL3qfAIt97EeTjFyNIm/Vh6dmc4UMtfr+6+OwCrzszs9
+0YnnvhTSdZHsr049IY4SDpgG4o34ZA5tIA6QVwpx8DY+e1NtRsR18ezl8+gSJIDR05qAY95ayte
37wTQiwCPcj61iYqGl7Z6n9sHlXI4GGeEZY3ljOJw7MmTWNtkjU9ZtW0H2nk0D1UgOC8Fv/wU851
ybU23cJkSCDAk/0KFLnP3e2NgEmrRl+TrpZTCHUhYg8byb/Kgr09BeV0iek0i/85zwrSRIAt17b9
ulZg2sSKgAHDx4fIMc2EeUL9ln/hDgr84EXIDivAXFEBtb8nQhqI9Tr5wNl3sD3pNijFyWEDdAX+
GpLaFRQ4CJ6wri6DpmnM9uJPLZ4ornsSqRNgzU1tapWVxqNUaYhaR3M/UVebpPIvJfm9yqtYH7N0
jfPzPdfxtgEkE/rv2Am1QDTC2Sqv/OldGHyOMQ0n/GdXzcCSOgHL9iz9D/PhnK5DQWmvUWPkffUa
XdfLHNXx+97gjHswi60V9yqkw3lITSGmVVxzHC9h5c0cO1diLnSPmeHBotDJH+vEI5GVreTxTfNP
tgmnVDXnjZO9uiqG2opYcahQ/ZDwxipjdJIydJAs7RsZren6Llg9aQRI2h+CVut2QwjehTfHqzRK
srPd0ruMm99t51ZBjehLln3fPF7ryVEQsrzCBdHl0BJSVpQMTHl/D7zycrG7yqvTjT2H5lgazFqV
PfMYVanyQuN4lQ5Oyv5579mJ32krBnoQHwtZuE9Z5Vk1mm12jJIzXLkLqJiA4hJYU3SQj6LXW2XM
CWDPCfFqeMqIGx75ZjYZ+m7m5/7Tqf8AxftuxnX33F3Lw9KqBn6nrwFq+LE6Q4TpF6mEabUvjQTi
YARhwTuRJj2XRlniNZlLyYIPD+N5VUf8IgJ04in8boQq/yKTi8Mlqgj2p2OhebK8FetJ0abtj9sl
Ee8uS9J8oSMvSnfDMRouVHKFmd8xfoRFvxuVxpcqXfwy0fcYMhgmIw0TkVkl4BG51vDqO+dbKzH3
ry18QdcjFAHt2YNj2PMPJU9NxixAK+csXqYVWxXBe3ZkeVTu20V4a1gMpUhM2hw6T4LdfS5dWZ4p
54uNN8Hip93gt213lOn3L5uOyAaNyBHhbwNad+wd3ybJ5AkykVvdtsmkwt5bidIKs0Fz/n4h5I8n
3u9xW6Rv4fcBqDHKNJjx9yeuU6bx7HTrcRiy9D7LfcPQCTY0l/XHfaFjAamVAxeJvtLRu1ggK1/9
uPF9EVdtyj9h7I13mQL/T34NVopLiapqTTdCsXl3nKNj6ef1rrdx1QFqcV6lj0bco9ns2rrqoASn
Q6hqWx6lyZVxY0FRbLJS5ylaxZCi/I0ikGCg2Ff0RJI6VFyANi/4VFNRkeHfEdQzChZaST5AIZhm
XvJMjP6GdNpV2w/Xo9k1K+SuDAem6GoyJqMf01ycG4kzTXJqjIpvz1OHZzUoXQ9FVjafOFWRvI3D
oNbd9CT+TNY2igWjbqlBU+7WsqpZqbSOIBHmypc4wDDfXWNRqUwOnhegmFeHva8m5dsewPjDYHtu
+YuVJrXubZbTIxSrL+nWf3/bkZZc3aWPb+PS10lNaAUO61CoFW5URluEaLTTNZUYD08FqMscJYBa
nuF9blnq7oSYD3nWDKuayHi0Qi4keaZJqhDkyI7k4hfQ06llfQx4qAETDFPLEUl8X7oaKTGuMYwY
XUMNiUiUBIv8ZJLSy20LkJ+6ECm6ZAoR8dRqKYeDwNzK4wmqGKPhS7AyxH8sgdf/pXKGjNj9T1VS
gWM155d64K/WUfH9Up4O4sIwerMyDI5+Wud4tZWjGOFaVcqEaBmZYT2af5bR7nnUuDktbADbx56j
S/FWNNYVXK4cAxhBED3DBEam6bhCHqQT9OUkvizkkX4Usq950GPMPj6NAPh9WZ5hXv8p0ut7l//N
b+DLdZ3Qp+33iSOOPTVaE+F0Oab1Q4wNUho6lt4qwlexfU1E3sfOXoPExDRtbQigzKtTmyBNVWUv
pR4KIHaThFXi6Nt1OQqHH//ekFqR+CkmkxjUcXeGypIjy15LfXAoAq9YoMnCQdr2yh0mNjtNhU0N
cfRHSSSSzNYy5V6284qDayksiMNtSfcJS1JRfuKlSCIrTt46jBdZkbAg94XStUpuNHPHIexPDd6H
3ZNpHvPq2zLPVYDmdYQYHUASiO7GbGWszxBYQQLDqomJu4KAQrA9owvMDsqjVkJquj0rqOqYQ0ph
004CKnJn/NTCBu86xzLZOQMoJjmOitYWef0BZkEPClCw7kRIc6E9n77IWSw4J4+TNpDRMqUdCI7R
47a193eESzME1L7E2a9uYCjtTPnOrzDrIfdNSbyCSGjhr29yHJA6kvTHxVeqg54N+um1a+/eC8vV
LnPF7X8zR9tvFRuxRAy4oJvImEO4Zm3ehjD3hFgynYA+C6mharDGQmuazkpAtUJbEXszyFFxVwWW
Lw68Kq55MiaZCoO0Bh2X8n977MDYQwFAH0gfV8d7aExpaCsb+8K8yIGezwJ4dKeQnvEcK5htV4Rj
s1hIkILJoqsvHbP3K6eIH3pjTJDA/tV+iYgSPMdZhfeU9l2ZH+W+jcnNDsalIdIoKsQZHx85PhiY
e3OH4odBCdFVuN9iH37Y5AHtrhMO5pdYtGv3WFd8n8YEDcilgww/F9X9cv8GZv6O+rfqHf1eaDbJ
duk5fiyDMrgdyBsiPWLeeA/6PDJI4CsJExBS/asRfLjiFTi2FIW57cNGt18BmL+R7YfopWJjB6Bw
SoBxEh5jvEd0rGmND9cp3PyRrrroT3K8aKmRi8cCZWNP6Ows3hskjjT/a80uiyl3S8HzSGEJIKng
+SWb8N4ewA+KCo29sZ2rYMGhIuRpUOmML+Cx+fZyXhXhlSnR0ua9XFpaWbCgQKTTlpscbMaJbNGo
6Rsa8fn+ofuMuPWH37283Unmf4nCxd2F6AXRlAo1BR3NrPH+cK91GvyuodS6Ivfa38/UuhV+kPYf
xujGFwgA3qBnt+gvqEZJq69ZZjIDWcMYpcFWRtsjvpCdWYKBNG+M5yLWr8/4Km4AuPNw71EKL7yT
eMK3S8MkJWQ6USU0FkV7y/rym28tH40jx9LnC1trubHMcc3O6zkzWHmo6gkUI0XJeQ9xN+cIIAav
7j/4ul6Lmv2MNoV1RuDVbalZNkWQNeehxhs3pdXy6CJcBLc/jYYbBLNfo4L/D+JeOdunOjq6/Z/i
o8D3O7vExbkU7qRN1jX+BIxJh9ZJ1aFDRGO7VzzJGkAUcHBgF3CyGWVmXkP/aulyY6qMdHTTrKYF
KskJklJqVVebSHa+Wp7H7l5b7UrbWDSAuw4ClixdDnrnKaqiyzdRuf+R8saqN60SY9xIElAvKuV0
CMg8sTSWohCwr1K3HO7gex3MDXp7cy6MzI3/u23lVNu//CidfedQURByqZ7Y8rJXCnuzgCIDOCNP
9dJpKvfEXyQD5k2zGua1XNKsqbr8kIrV3JvQW6nfNFtkpgjaAFtdD3rGM/1ro1b8VnAI2gWJ7Egx
nV9+9WE+a4vlUvr5nJubwy0AQpJwHujCS8ln6N30rCl+BTWiFZuostbAeiSrAdirN74UzUDhs5ue
ZLatjJepIoccS9zEN2YLlkJToTLvdAKfGOou8Rl26mOA6ReEcr8XfaI1aG64bBCZOU9XVV0hfvmY
3V5YfJFdj1P6A0mBe4/Lsfn3omfeQ7P0u55W1kdRdbke7vC18NcMrvvAkXIG4FcXVaX9WSFLvsMn
/jEBimQ5wQRxDffNweGgBAQ5/aLxqSH795GMJBP5DFWVjK4FfCB9uJ1qaNgEa2XUmonT16+N5Ce3
9YlMKFHg5yYKCXBm83ZHzib9nRMQgWIi7jJ5gklhMdmcqSdTye7WQXBbfboP38nvRt0E47y3lvj1
5yjADZXUO7v1RP6URbZr/ZqiGDZp/74K8lJEwW8NqfbFtX90wh12qvOZ2SPBeH57e17/ZVhkTwuy
ipoz6zhl4t/4vPopZvqBbhtF1UsZKE3/JxJfhpEJpyfk2uYSLCXN1Qz076EQBffz6SwvuxIkTXU3
rQDFMcw9lBeRxW8s1vZMImdekSjPIvOXMp01s0j/Pm88S/OFhynRvU9rrlUGMtdvlwT50ep7l0vz
v4I/lKHtvPC9uStJQdiE2Kuzj87bX8XL9puI9ToK/60UIJIwBkWEBl+AeOIZQuu5ZoNZFryc29S5
uOwB4IbfLgh37x40OyRE9Sv9ZhvHgaGN2TWYIXLtJSo9DyTfaLk6ufuq8c603/aYLhqxlrAeK/Z8
O2dpZTTFerSgzr5PjbzOfwUD0r9YFCJA8tUQ0s3RKKVYGuy5dThU5BGz+76y9vMVbJUhe9TD6JhL
rePICZzMYHJNIMKNzbEiKL9wUeI0Zt2EuFEEebQllE+v/m5keVNdFkmHhbZJTze065F8tcrdjxnm
0FwHqPcmMgzzb7D3r7D9EH94DpLGUQGRZgIWr5CX3hb1Wvf88HtmuNXgKhOLpWcwiJUffi8eFvjw
zUk1J5VcYVO4udxPIw3tLGZGsMQPkpJ7C7B29T4ezmTBzu1Y0d8qDxbCkSJdvzqjri4tYAZ46orY
9rvIHoZ7k7+EUq1S4y5W8vYHfLRRu9CBmYIrsguVFrI32+haCoU8XOk7kwA/8QmW3hbyAMaJxvQ4
3U6iZAaCajl4t5TKEBF2E0+qh5EQfezu+m+ItcHNfPzxGbbxxtNYupWPazqqOkJXj8rJ+qhKgqmx
BnpYsKg/aVahRX5fSL4XmzMYn39mLcz2Tos3VAp0IiRQ5m9WzLs+jqlSt6d7HLm6CF8/8bD2+brj
PQwcHiQC45qQxLz3KqdstailQjac5biZfVP4McPK+uTVW+nYfUfRyEJy0zHN3rxNS0blZH648gqT
0qZ4dwbkGPoHq5xd3w5qUf9vfAN+XjSiUkLLtYqzR7wB00ZWpKSmnlbCSWzezyxe/lxrOzsnIElu
9bB4J3370dDts3//379cDiJNa6baACWtqcKlG/ftHfxhuLBVAAyheRApdQ9OEZv8spk8jvsqV+aF
qWHYkgutEIQM86X9AGRyjY62DjYCDK2Q5bN4tAAzDMylpGgEt/o0DCfIwApngaFwCait/e5scjyj
0k8NZWzn/ss4LAuWrdU9RpnD4LmgOe0Daaav9p5RqbK2jHF+lmM7PP06uxiHci7vbi34Fnb0ZKO6
4XoCzTHKVnyz60tJPnW8NptZUPnbRvAtCqyLcti8XWuVBCwizKvb38ZcvCoR5IBOa7TMt/KI0QO5
85HN+5mgW78gfrsf3gnf+FLgUC1RpuVjkroFAnGXIH2oF5bTXgYPqB0YQT9MWImLNWEpizwBsZ39
vZv0zJS9yZsWZ60DMuPZyecgFf+AFRBWShkK
`pragma protect end_protected
