-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
vgTg3+ynqA3kUPKKBmh3wWWNJpDdFxnp92vpwlGD4kUmOp6rJae9X1fa/SBpMRAW
oLmjSRA6uUQTEa5a5p4ueibJfI8wxKQA4xFfAiC8vb4U7l+wLe37LbrTKPC7uk9e
71sEdyN25XKprEbVQokY9COJlSQoF8VowsiDJ01gF3KCWtwlkNRyPg==
--pragma protect end_key_block
--pragma protect digest_block
u0bu3GDF5OoDQqBXv9OTCC6iaXs=
--pragma protect end_digest_block
--pragma protect data_block
M0P0lzNKYu+PGK/q+HLaTDyKlAC65ndIeQWLEavSoHRfI+5/UZtKBuTnOPvca1ko
tXbCYhCfqfWgp5pMhpS3gG647Mn/rvoSksiVq/N4wdXHzOj/tRXv/O0UP/c7+lZr
QK1S6GWCvws5OMMeLOZ3jWVr1iraBlHjsKIE/ptBVxI8gX2d/NE2LsrmQaw7Zji6
bTf8bG0vQd33uC5MLD4fR5CYrE1xYbNW6+uERGy7aglDO2S+c3BYWP5snFVWcXFj
JMIj0UQRKE14jDbBmKeN99CTJRQ0nVeC8hA1toJuar/vsTjwqjhoD7PxRGCr36UO
uRobakeF1UdW+W7+DnXg0k3a7eH97tKYFBXE6ibvMwhooUO5EJKHfTSoBtNQuVK6
r+WS7o2/bkUirhW4hEsQt/s/laIp+gGKdiUsMYj0d+A0FIoNxC2IWHUL3ajbLAO4
oFbPpX7/Y2h82EYfEfaPjrG6h8sjPIg+TVSWnlYcENRyAN6agn+QQTZ8Us6fuhfn
1s6MhfPvd7w9g7Qv9ZrIfhk5ZreElFKb1MYJX6CUXdCUCj7Z3NmL9Ae6g57j+skF
ytJg2dZvIb4vkwDywcYH84NrQwn/VDXFDQgF4B7Fs7VVeMhhRJBl6ZHu/FrXt9yA
urQTaJVgBCBFzZ68vOMZT92EUxBehDQO3zDZjBc+jpf4EBD0XSoN71EGtjAyE1SS
yeWJmokvVxucHkQkhboaugc7GRCBZ/tWjVdHt9DmuLseRstVZm41NYmahMn6BVgk
zOToChtPZ2tb3xoBkd/awFOluDTwze8czHHpmKbBDTc33vwDxkib/o61L5De149A
t3aDC6nK7uaPsdeIgntB9iNwBlUaIENSn/3GohrQt166jFVWQ2+UdVIL++rGXqMp
n13q59bWFurW4vqTm53GI2OUt+A54tpnCI8YEAxF8cirEqSS/Qseh7Oji8myASEK
lE2X9jUzHF3spcjNPY0BXEPN6Twfue/BjBQHilrHMYIfFDk4T/lPOKpPwlk4zD5S
OA3FL/3RdtXkiPSjhuXKcWTbLuLPd0ihsZPgA1P99J5O1YNjCGogMUn+x7MJE15J
1dOFz+fI7OUpDXsqyfKA4C7TygZOC8OlzdJvByRz4VpX5BdNh5xAPEu+Tgkh57No
Crvl68BnCJzaE6sxFVilJM955WACzZ2NeDXqQY+9aLN0Qgdl9Y4w8A19vUCjVSfM
E0ROmhf+9yGvJp2gpsvE60Rm//bwuVxIsqOxbNQILWGaPbHb+5lhgXNH2U5khSv9
QpLQF9YapaUirTZX10+aqS3X2hSQNv4N8WtIRx92GAM9BaAn+rsdVxyMatZfQytE
2tJla1WBsZlwcW1MQfG12wQenxMAnqXC1OjMHODrYXjI4svXdwTCb9blUgHP1XsX
uf0SFlWBH7KcIor2AmvA1Dpvby8eAJ+hMH0g6EUNJDSenOxXQJeKuGWerMKIcecC
gsh8SEBNjJ5/TwSzRi8dC6kmHMHY5OFzE8601ZU+rAqX41rUKxGfzSPp4PLj/07V
UQ9AAW23QFy5wB3ASTD4pFb4aPpmjFb74hDQuXkr/zCd//VlXNUK/hDrJQE8+3ZF
deKRckI2MRMO0zEjZIWCwcfD/Q9itWWWp0/2pq20nISvyKDTBxZqf2ec7NguOjr9
VoGf+PFzcYteG83e1gxQf1pHkgdxekO6XEkcMjHObbau3gAiZSlZvk9nCzHVc4at
7VABWdktQoF9f/cksaf6EYUrXmds+QpGZVBJRLO5h+SuolcidwmVRY3M7dcX9kWB
3flt1SuyjQPJQ81qlRfKSO7SnfP1asR56GKlRIwwQ6v1kqFWDQy31xEI8qo1wRLh
oHHy/7AbjlXIjB1mOzl9vb++Lq1uq3YzVHtD+WVC3pvl/i7Ahd9jWKpeWHUs7gsb
tlM0SXfYQkXQOG2HZQumX1wqKhbUr8uVxxnWDsyhqxz+HNMDrrAINwo/U2rdcbGG
nLZey2NDcUQ8IR6SaNngKB1qxSqD7myNJiqJLnOxTDEpePM4HAhlCSuN+9efYYGk
2cShqtIlg0QvPOzhckl+Pp3xtHPJxneghBESHC1yr7+Qm9BcUklU4VTrx2z8IfFt
qNqS98gBYLfEma/TpIxTkYdkQGZAcrAhFDyoL6SVE9Fq5bedq75GRIXc3KF8BbQ2
ptFxel3TIewKjB8q/NnbqVHw0DgmfjlNM1eycGgr1gvF+0w95vEyJPWOOYzMTQeA
eJ9i6ki2fTMQ62lkw++n9iUVTEQVa3l1sD6RjZlN1L46XUB8xqrbwaG31d0CQN+x
M4iplkDGsdgQAdf3+tgyMiuwQ1H41J44faOK3XCB+Mn2ya4Ub8W7WoRFlFJe8Ah3
miu8slQhfLVH/jTYBANX2YYMrFIpmtk+CoDPWmxcbXZ6RF/VphiQY2sNUYeARBAp
fPG+EACLXvAalwh2i8vrUoFXAyZhw2hB7akcz/0aK3u+Er9BhmkuYf3pwG+Rx58h
uspfpi/zqylHD9X5dH47O1A30Y+sqYra3CPfYo1OrMswn/K/BJSQQMrn9eyArjqz
56X+VHopYmUG6ENrORB1Eyw31wrLVeA+lKDTuQThmVcux8ossB1G/mxv7fLdI2q4
qcHtdWunV6TFgDJ0Y/UW+TXnaDG1ovLYmqf9R2HDjVNdGbMlzn97tOTu1jU/ly72
KIj6FeMclyY27eNzKaqSDUFn/1tDo/SjFIIDj/54JyGGJV5AMj9tO9e54eQSzTv9
/spSJv7SmAJQcvJsyk6gtJ5CPjs3n8BoDD7qMI5lK2wbc1H9brorEn3MK5igWjFT
xVupu6L3Wn0UMCEjbUZ7Y+1me80WVd/7cSA6K4jJTlrzJBcKCRpgwficQXAK1C32
N7LpuZbnSWoFLMzsfB15tP0wY+Xq01KCKGKatnCeaeld+uMoqtwCBw10J4lE0VT7
1JIaDo9VZYcrlkXSIqF6a/TbimVhbkwsecEHWhqSHR2xuTdCJBwWq9mp4mi2685p
+NJVpYy8TJpI4dOxBF3HHboyx4cynCss7OTmEA1ug9mBgkEr2JFvRcxmzorXjWNy
Gn3m83dQGdM7bojaf2j36hHQOhBHS83+5AGH+ZJTSj7B1LZwnfIFrXghfwfra2ye
mUbZxlipsE9vYXXR1I8Z778kOiEtNeFfd9SPdhR+YPrMmuk9pqZ9AbNHyImeFpV7
/vo+yCxw48UU4wpYSqFw0gems7sbyI/wAx7HuwHHA2eiRaF8jWG9MsOif++NGT9M
TDw16BRYfL6neh14AkdY9vYJSrXPaTx1tupq1Z2e4ecVsRFp3utsb1dpJ0vShmon
SjJFa8ZO2tMRgIwhT4hVVs5OCAIh2oRt6nd6dlAzFm0UTn7lElxoH4m1BSaRnzFQ
kXfzIQIYwcF7sNvyGXe8IG3FuOXjqBXBn8WG33DLRIULxThhZ5Gq/58eSV71k35Q
Cj5AObMgpseIHLHe3f/jOLQ37wISOfiWeDOx/DhDGSL54GeEYt7Uptg6tVXiRj+a
D+dDDSUTUJw1MdZllVn997/ACxbOM2GcucyyY10iJoYMVUkCacnvfUNLm3DDAZ6Y
kdZZ9gaionjIA01LVWrFPloncdMCOX9aJPKQ2xnPFpi9hqj8p/InBbFMjRhkMDMW
Qj4CxTyB+tP/x0CGaLAxxMLn2hM7p4zTPZ6id9d5MvyVGi+cfoIz3HmxN9GGLWzA
DbF/US+numMk8Iey5ynpep46IvTXRHqY60quprED8quvd/Iku+N+bBnzvStUIhMA
DaDk4iIi4L6NFhzN9YXpWw2YLMCaLZyq+thb+yviOwNmwFmi5XouMvOqIdJ+MACL
Ednrt9lFxWOgBi8IrXVPvaQe5babmYQDi8emUwRPVXxWtJQAbDRaAuwsSi0qSQeM
MvJriVTuT5DyRuxjXMLWM3zx3R/liKs87/ofTu0zLegyTYxwr+fKk5cWiAJq7xW4
c9yydOxDya7t7D4puHv6SoOxug9QIByClAMHv+5s5PKAdK+ac9t/dz+iQ88xxvtU
bFMAp5dSP2nBRZ3fF9QRPKwKv5kqEZsFAp0by1cI+3p85dZqyzOQXStE9eu9D3g4
w6GMtn4VmaWfpuF7ARPLpLBcmdS3R1rpP6tml7iHltEY1sQ5qCuO32blFKHeDALI
yo7veaU6o6lmlfUnxXsJYwpK+7Awb2RN6yvDamteuvKuxTD8w280IKUqDnCGCbL0
W1qxjBTNZXV6dJhI8Ey2Ok5kES+vhhbKhpTD3BZazKYWIN2OxshXSkdpFupSmGXU
vOPPnlUIl+UtycpFa8nWYuZycXrzdneoo6HIUaQcOkBkECf8Sge+1tMuxqY/MBQ8
Vg+yzxNc7dko6up+AdkCfIEzG5HXhXAnISGOQdYctCo8ukM4qjcEnxV9yKv8ozZm
vQOsrjNbw1gsM28Kb72T72Roe3rWQzvX1U02KY6Eqhw6H3mIhea6ANN2cCKAjLht
eyXJzTfOlDcU1LLzia4oI9QINtSigikTsk9QQfYzz1xBiYozSgr4GlZ7Q31gOXQK
jzRJ9EZVMsKKSFjvPr3x8XHTuRRZS1t8Rj97h8ICZX7FLHdG/RCnRFHmaq/N0F6P
sZtn/eZhnTJvzsVdlZjktHCsE+gthegY4FYOw9gk/fO3MMO1hW45avsnYr3U/qKg
8d7lflj/HIsVIJfromQHWZxnH7IcAnkJLpXT96LI1oi8hWf8S/74JVUkB+19Nva2
GTiUxK/pJUSkhb+lMw22dALawKv9VGIrSNHCztkoLh1dF2PFol2MPB8xc+EE5c88
gCnpb3zY05VjZ6WcmtUm3q/bcxRSH6gTui2MScqUssVzhWVxr9xmM01vSQRKetBn
GqgOrMzdEDTk4XjY/4ASVYhSe8o/h1nbBJefEqtnGLaBtT9VSv3iXKRKIeyI/VWk
pOFnd4o+TQIaiKnFNKR1UxrB15KtiHfGm4e1cfG87vnATJT8v4eJ/ROfeGUrUnyj
/6OOBxe5nB+lJIA5WlwPYh1padg6ZD0ZrHbGnqPm7L9T5c9bolN4rAYv4VS1ek6Y
vAUjqyoaDPXkPvUcfRvFu/N9TFN7nUT1cO7MZeCJ9+M7zrAm1Qpl/yYhi6QS42/o
/JRGvq9uqZflhTsXB/natTs8GUN6/WK5hGESnTFsSJrohnVNm4wF7fd78wlDAL0c
77Wpl+YKGPMfiSmn9VTBSUeh1Nur7RvfvqLw5zCXa23rQyUknkanZ/ZirFSQ+t1x
wl1UVjvt69tfd/6Dp/brapLOoJE9u0UTpIGgDDRB1Cp8fv/VfCMMBzmIJwBHAcqZ
4hDmOrLl5cUmX/DvFsj18mAewcuaXNzgQsBCKufgP1jNUYCDCydJ69tKgAyHUFyl
rpMFxV1eqzNpcjIxH0+YIomkvXURCfSyp408mS09kyaroDuhITkMITQipndEWZS3
LbUePrNUYy3WYnPBFoaMwoAVHpvHWxnnR+Hv+yBZtg5QCMvHJfObBrH8o7tPcBu+
wRHqc8AEvhVQf7tv/FmRk2qAL0rSnV/8dyW2YAmaCHb9YP/E6gXPPX4JO0u+OuZm
jDxOhb2Bp9Wdm8Vh9uJ2LWgKdX0wudv3+4la5urBFZ8nIurTB/afQ7nDsGGA/LFH
lCbBFZ5Lqlarv76+jq4/t8XIPdPn1K30IhBqwI2RdM5/WL5Ly3bYKY/ywlXUVS06
G8bk8S7Q+BZiloNAB22vODxIBvBf9lywM2ec6reudHcNiViaTH018oDAJ3W3h72y
QtUh1JEesIUkhZTKFpeAulASwq61lswaTtkS7j9l8ru5y4HZyL78c3aa8lTisji+
/Zgcxe9k+bENtgGv8F6Xfi6gof/ZF9m5OSI+rmIHP0su9ETiMtMILS+UNCUD8+i1
fHdx8h2KDZz3JPOxDPWbZgzK/RTB5goPcWUPSIziUBKka1b2nf4TIq3iisIzb2y5
LaYPFNlYSw0iwqllJPcxD67QpPfU78V52xlvPSRJcGDzE426xQ9372Qg/Mqs6anK
GMVYLjRZ5kJczhTel0zZip7YwTllsJxDff5d1qCyzhbP08s+PvSkZoB+f4ag4usm
nRl8mUu6PJmdczE5/YZRaiDHuJ7tBxvsylAxDylIrnQj9ZDO3OVbwjW5hDuuUVKm
yaFK6nw13cur5sZfKTcPd7ikVXPQVXw5dk9+uUafZE0eDubkcf8PPAuZ7ePLBCDI
Y1vloyEllzoVkgUfFHzDGSji9u5ukxNC8bH0nPGaEaKkkUuJNnziTpNXg+8UoKEd
bLSlUafRiebQyaxVH2R2rGmspmHhzIMwLeVeRNi1JEQFlhY2NPvAHPKx3J1ID1vu
0cCgvNPHYNLoU5/ruOe0X3ZSxWgAHJFKSKKiYYC4634E/EtuzU/wybu5yIAzJ4TX
bUVdJwrM3kSt6yKyGvIsOduZi/oVDG9Weec5PkOef04S/PZRtHENTT9nYLwgbSlY
iv1Eick5iVLKm1uqCb/81S8N/bBRObRtfhuipZom/VS0dGeaLY+TTHXxBppZHXaq
KUeJ7u7P49p5/zeG2OI/lXoXujsGoSS2ucEExxFAhXWr/Ji/xUnYBKp5bnInygrS
AdxDiSlx6EsKGILOOGLdmxEN/U5skwa2P0tQWYXZC2XI2AdTpBtXA6xPbTGvnL21
5J1vHqes6SwuNzKZYriorbNekDfgjegchiaDdE0w8q+WOWJ0zI9VVbr6k8LmSYgx
ueFFBiOMIaDub+TRnxMHmevmQ3s5MG7YVkepN3qHbayu5EdCuJazTqWkjuY7xs4g
+LS2BjCcex1gN3nMQ9bWdfjFBdShmm0lAADoETOKao5uUhXRy2Kc7fpIs9dk5nEc
N6UvzEqVLIOaEyGK/gBbPVMUyfRUZABMIAjlfjkzm2+wCrokb2HcmJvdrabQRZO7
CUZxPL49+hD+BBNenSxUlOrMiJSE3sisgCWZXSOyzW/sFJ3O5eitthZqkB5L6Cf0
E6C9FIGcpuybxUBhpOOUNLYYVwmFIu4hm8iz6oVTAwUkg3O7xLucUwLhi1GxOC7E
Xq1MuTnvL58xDZz2mcOM6PJOs084p8bdiT+eLWLZiy9wzI/+ljn2WCQT5Ad5Oy7h
YNZQEGm5Dn2YbLzrsDEZ3v4XRYUBCrOGXBoxBvRw2DUou4ueirzklH3pIiUWUoB5
w5zqCe73Y33BZTLNRtjZhgO/hSMSl/D2V7Ke8h6bc7eigyAl1GWk8gtjEfMcivhn
1rvlt4xTExqCpZ9KztdI/ua1Etrm6ZpEUa48NsR+GOdxH7C/ThvUGl3jkX5hcZ2Y
wZ8s4M7UOxceccKSCQAuG8bjlEK0y2f2P1K0eQpb98as75QYQgXtbsnCwN5RptGN
SQBJ9iUK4VLgSPqnfgmoFaG5a78qCIl8btfXgNM3Ftk+6P5LDwShhMHuFVpcBteq
2Yzpzv5deP45WjWspw4ieFJ3XdaWwFBiPgERNm1nYQ0q+fqH+wSI5cXUitBRrRrd
5K32iyPj0TwW4RigYEbhtIjW6rclwGc2ByNhkA+a8QibyVMbONarWmoQlg4Xrkxp
FwqZzKipgbLDXSadA8wVimTuvR0Eq+hAF7SbHtrAfZr2JYooJUd1k1R41jHdKg3q
9njpcvIKHfKoUFOB29nreQcNkqRPx4pHjo396zr2uFNZr69GlQD8S4c7BLQyvwJl
Sq7QdbSeKk6lrKORlkaFPlif1ld/Jt5tb7gp7az66QgmtuFw1kHLLh6xFPllmJRK
PriPtT+nZnLW7QxOPLtyx3Z/bUBd+hGAgeGHZq1SnWeX+Q91x/N27aAbiL1C9O16
4eRFCZ+wPJJHVGTs0WyJCR+0dscxtX9mHz6/bdbITOoh5Zq7RxOV/mZXLtFzuCGE
0nR58KozXmp1ZMC6ZuPbBTtnpK98uG7ZCkKK73w5LQq1zdDuBlsaepIwvlPO5gbD
ezLOOfbpreXSTNyBC/saIPmeCAxU+mnVpVVJ2Irbwi+Prw/Rbqq6d86R36Y4hJqn
tMGDJuNUvWZGoEuFU+UP0hLAJw0ttfZcN26ybEeNRzW1WAXWBhnDdITKp9tozvQx
ezeB1q+b6zEVqon4Z6/Z+daSc+0QuxO30ZIuwFxVK022t1L2EVsRrnCRq8K8cqTP
Uj+TNAZ+JFx1GAjEoKRGYBXBceYfrT3WelmYeHT7a5t3LD8dvBFez1w2rdOQ55Dw
fdVZH8Ce9JvYdRpPFFtrFUPj6A5i6ZU0pWWlbkMzGgIlQyoJUR2WmEkT+3sSmw0x
oAeUsnvdXPokCuKdtcpe9o+P0OtnPe6zpJNk+RTYEBC70EQCVL4nfQvqYlSwhD8D
Bg5t+V832LU12ewqL9c1ofIGyYbBHmUa32Si7tkgDK+KGE+gKAKUuieilXIjG0Uq
v/L26R7ORK4Zezhomvk4TzlGfXxBs6phZb0PLb+sfFSJPcmVM/s24WJUbAnKrTmQ
XEH/tvXvPU9imzT3Fr+bM7+ElBRYxgOLZYV9rVHQ8NMJNr2huMpgI7uwphrrNgBY
buu9ns3AGHbCfo484Cq9HA8+ehN/Q2kgDmIp7YQJPexf83+Xe1sHLXvNiYSaQirG
KJvSjl5uvxwA3ykydMjMLF1XrHBdHuZvY5HuWEp2zMhYxl9hetKfN35Mt2/O1N6A
m8h406sFJkSoFN8rbkUeuG8+PS3EfT2W9FiCyTFTheWSiTmLjfmHgi8qR1xn6lE6
SAHtEdcDec98T6XEUgLfeHhX3mvWkRLqUFQm5vNHa2Cxa1ZhjFAJdzZoMhZW0wHT
UIQQHmlkZwpytMEmIdmM3kbN6C0qU5CzsF04F1vOXKk1HhJNixZ/H7GF0pi48STN
aZ335uEo6EkAteNF8Mf3oXIaxWqBnvOw4/lBN6VKyCk/QUjYd2knI50MuWOSChPg
Tmv6DcydwiA0pkjjf3Bbv2i/U4J23WcNvPYGjjmyGSxCZfQNlM4Hiw7sestAksZS
kwwJsYbtj1aqLb/O3gHNjg==
--pragma protect end_data_block
--pragma protect digest_block
NRchKoP25EKfADAvzSAeanz5hcA=
--pragma protect end_digest_block
--pragma protect end_protected
