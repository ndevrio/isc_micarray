-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
v1B9LC0jv8D37bRlEI6OgZ+ExdfyxTyoPJDLj94ftyC5NWKgK3O6i/eDqk0MxCMoB4ksKW3CPRZw
1kFg9tvWpGFfLQb3Qw9yAJK7qdUCplXQzM+lvlPqSlU1ie1MF5lwt9crTLddcwl6yCnVf7Da7wsj
gr4bTiBKbESRrjlJMpYwbDyLTLK9SCCcjB+uL/M8LaeWY10B1RKTl07sXcdyJ6gnIZknffIsmGot
x6sZ9dBAJxPm2pD+Rn58GEemn7DJaoD1DxG64lBA16UmWmcvObn0DiqAbbeoF2GDoeNgKBL7ttvZ
4xJdvJlYIa64ew7SmJCnDgGB+4TtgmlMN1z/9g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5088)
`protect data_block
oD8AJGfpcMwNqS/7nYK/cszpOT0Bt54uNs46plKnEOcjhYEUHe7thfDVhDpVmXKnJ2i279CHOM+b
LyDvkdvcluZORKjuD01aHcTKE6phI56kpaIwb92ukvFFvdlZGh7ossPKO+jM97E2SEIUHysRJZWS
54z03eVbCNMWG1qXfIx8tlGWFNfgtEP+de5hIn99Y7YMoSJxiiEg2HZtWqoVE90B1HEQcVHwAYgc
l5kJG4BmaxOq4Bsq7xjO1iqb+XkxHU/aT2/thnkWR3cdHL7ky9H3a5Bz6jak/tU3ZcNLRTKp/wx3
yGrEshrBHJNumscI268qCwxpsMllXg/csGDee3IsLL7B92Ly3s8O9yUEB6VGzS7ak+xq/cTF5pr8
NJmbg234KglO2qvlIyQN75nDy/vooJYo+mrbQtwU4K83fO1YQSmRKcM0v8ltPXzo8MGQZrdc0pZs
F2MaG2eumFHZQofLe+o0itKC/oktgVLOpRip78TqsWQH6LQmEyUKcarhI6/QmHae/30Wy13Qkvpu
Liwyzp/W4zmCz7aINwEIb0fdQT7xUmRACcKjvmf0Ys2r21oaBBFKxV5rONdFoj5mki1DKOI+IYrj
nhjLf/i1Hjph2dITFq7tCviQysa1lSLM33F8c/CCmLcludf15SWMdLIHp+6Vkx/Uwg8LuNcf62GQ
FgnqZwbrQWQTqA3LS2GVor8sUcW+7yAwrHRiKfBjSxZCZ9GGmVTbnDxwoUrsHRwZiQaIAppjB+X3
6vCaIJwHp5GX6SWicyYDhIv0596UDWqRzpJOxt8w7TpohlUCNPlK0hQVW+8Y2JqUoVDhYNaLabfh
XE1nIMcuV64d+fKaYqSwyt14XbcaOTEAndicbKvSA9+s+fX1zI7kFQpyyWeATGmaFXYCE/0MGR19
CX7SYzv31vS/FN3IN6M7SVxr3X7EmDyJ3furPRpXouEzyAaqxpzXDrDeZi5t4pyIV8jlbygrXkGA
zpGg3deWc+9m9+7FmdRfZJ4y3JOCQ3B9DHf1QWnDHVYE/CXE0SlfhHtnq2ZQL7UP6UGMIguwspvH
t+xI2meyt1n/+H1yF452GrwQ5xJ1xUS0NP2XY1CchcuKEXvLp7XGM43TJdeY0QT+QAjS978P5wDf
x2CB4BqgiQksPkhZJA+LzvAc9pKhh9NgTBJhLTw71Mq0roz308+ZzZaRXXoE2OW9c38eN1PNHy5d
lQu3WYcMS4Vf+nfEMy3Rn2po+AXFrYqSnYDJN2woA8sA4LaptVD8sI+KDPS0dP5TPlSgVp1ag/Ph
888gpfGj7BkgyGyY5Dbe3VoIEyibYU8V+52h+nGMmNj8JEnWv33jZmdJHq9FxoEkdLR+tM2rhWED
76nQzr5YoYAuA38pNn+mgbVbfG/eue3uOvSB7CQ1kCzH8wQIWWGQj/obIQJWVp3O9KoIO2vd+X60
crUAlwSn2UYCWJY5m+PYjBQ6wcQYyeyEIT2BCY/yEt1pe2+N80mg0opikPYIOP1HK9IWKhZ3v0/E
bc7ZUCFUNYOUL+sySXMjsRxx7sOF9KiLForUYwiDJqQ+8NwblFJZl70aSbcJN0qFU6/t5atZ/5Aq
AfaT0AYz5/dAogldUpoYgDQN97zGGWB6QyeD4aAF3GqVuYiSZSnF+0Hsvv7M49C3mNU3BpVmjLjZ
fPaG610Dq1660nUKRZsyrotLb6QcZ/CHN3tkEBs2mk3ywjNCdYM/FEAHyMhu3uJvtTTfgzowzld3
kilhknKnpDHOay1oGA9UWSlr7trA6u0VRyzoN5p+sVbVWbd3vytPY/uaF7QlW5r37/iVP6lMhYBL
uRJGw/tW9ijYdGrABP2OrPYdQ8Y+wppZQ9h7nEFqHDuEItNv1D00Q6VgiK98DvQXeVtuo4D1+fqS
TXn9hffSQX45d7Q1zc9rvINNn8Y5luYkAuYKzV8xIPU1cyFeP7K+TcypTfL94V4D5IYUAi0ckkXu
J4DSZx4R+EoJ78XPL12b1u2pZPMk5FAvdiPQDC+iOsshxkrkz+dZA1KYSSNT6DM7uimOVsxldlzP
nyaOrL10Su+KPk+cwwD6zrVjOM1IMfzPZ/lBEQHjxYoQcldVXAcSwPrqAKkvi9MyThJx0ecAp16Q
q3z0KclgqR8Oe0zoV8/1B3f2EJxu7DEmXWuESQPEjpRXJUqrK4xdypRCZ9xOmdo0FhcM7S0qnks9
CGGEoh2sEEDGyEMebqDNirBQ2P4KWLinXBFWFbhbhblJLilJsL8oqMdADcgDL6DwdhnX7sdznMsu
5M5iH3tGZkbfLCyOtB8AGw/IsrQtYhHJM22ctxexMPsKHyqZx26aR4pVmd+GJS2qKhI3ZE8pAV8J
Srlyi75LPErcx2u82b5xE+VG86ZzcL7PhHpm8U6Qi1xpmLKJMI7m5eprNnkdgS6ogIe0OOVeHjuF
izlEsmRdMepqYJZqEMvQPP+hKRXt5KCvPCyKgOMd5S41dPeYRRyIWlV9AAoFMTyNXKVSF6XvM6B0
wdSIAkc/4SDR2gICLHXXJsvZkzKqNCQNVcgy7Vwir9z2kjmyeL+EP72zvNqx5YRbcUcHz4qVh3V9
Y8CH/TKMciSMtAOn3VrCUzj8SVybimtVBe/6lbENy2qDEw3TZI1L3NzkE1vGfDuIbhYuyM6TdlyN
hrCfA61V1ne7IIDFx8mnT1Ef8gPPrkusoB0wCxFHCPn+CKn7dz3jFD2z9OITcBuxgarRCYdVkBa+
/dg4DxgL707fd2R9ZKAxdi7kQKkpkw5WtOp19aVr/02tFx2mYixs6fLn1/jkWy7W9h9Bib/EmqSU
MCNOdP1sfeARDfnRdXL/y1N8/gXDcba4k8MyxhPxwSULJczjHMnINtGWB3Cjk2f/GKpiFifO4b7j
RA4YQRSa2xTadlNI48BnockhDjI7CFV0ueKLrQo6dMuYJp3q//2OdKgIfkxClejE/tIKJgGvVfdw
nwnl5uk5XPAs0etWwzdhxk6HF51BEJEXsHryK7hR8GRPzEPOYY0y2Ceqe8q76BMSugZ7+3d/+VLY
K8XVoocGYR8Sr26Xuv1P0yzLQdKQqH9C/eM5irnU9LKoP4iRfuIqbUj8f6+Cc7Ti/e5NOwVIl9SR
X9nhaDx4ibN1lY+Ver3O8cx1t9nZcAEpwvyEEyYxE/1vD5HAgnbmSkxIenBDFm973vP88iIqtALk
1RxYQbtHVU1N2u1AwNlTtHUnZewUHIbk+eRdcKAG0PA2R9/i9vgmi3ibFDyGPzaWh2D6XvUeM/dl
sWwBI2e3tpFO4OhfYObkPSJWOJVB38SjSbQjwNoYy80IqMoXqmwG4vNlF5qedAMtdbW4LXetHAVi
SUWeoW7J4UKyvgusmF7gMOx8V8R3Jr/nypzv/4UPAb6C559KXZt3eRaDE8KzhN5K1xTEes43ieRc
Rcf7P/By8ZueoyGlsBwX3giCuysk0Nay6nADpllgKCY4DMekFEzlOaLV5DHvc7HCAnb82z+V1Ql+
Chhu8CO3VBWaofFFw1+BYeA3sCdYaT+lLTHgqVtnqMe6I99j6XoLHmyhimyshP3psJ9QVqfHSCWL
ZvsB3vsVRR82twD2cqKnpjuAbiyqJRFGOxSBMmXsp40rXECIAT8x+Gp0jq1rZp9nLswIu8ocW3B3
VQZCTkJ5R7otnWDKVTkK/q3IcfRMxegZqTgD6OEAkBe1tOCOoo/7OXhhzATXX57IfP+nV1/GDUT+
0FYVTKjr1xI/Ki//5qnDE/CCnWgGB25u6huxWm9tvhIqhlgIuXnE15UulEVQiJBuCnkkaJ+c194Z
t6HrKzf4uFo84nFEwx4Z5GPVTCYJ20q3DJGrto0gK/e1PPBU6q6HKRqfmN5SuZeMkBqntGzxlM+r
kMR4U6akpcFJZqeFFdzSImJ+YNaMuvKTogWwCD52RKMMlatx13gMxI1+bm99Fz6ahPE+3KfYPWOM
aNc1XpiXssgez6+lVZ9Sb44PbzjQW0xHJSRWlApYBwt7PXbiGkcQZVfPRHM8L1oidfWOX2baLah9
PiXWwKST3ImMEn6MgMFCZJbz3xXKMsHkLzVlNBkD7IHWw+u7TaA7DNUq7efDAaU6zm27Sn4GjmAp
+N5+lBnUU3EtowMilMpTv5XCegH17669+Lq3FO4WZkbu+enETusKCp6+j0N1MRQuRqu9F+O3hGJQ
V1krunQdGhhnTQHPJzJfT8+ab1MkfDZnxLx+tt+X9WeZZzMW9s6kMBszDJbSYrquGnM1NgIX9aUp
oF/LSdo0DJim7B4F0N0/5KztSSxMqhECjieDy/Bz2zDBoksOWONdeb4u910RN7H3ez61dTC9M7Cz
2x+cgtW7zo4x+5ifB7FWST2iOc9fUVKvkLWDGpAi2FymXFxxPhuQ5wuPDU8f3p5JTOAjXnTELeyu
cg5DCva+AbjdSsAI0dM+ufQphOFbutjitpP7nn0J/0yGGwH0KCvkEm/I2uU7SvsB9kJV3JPgxZ4h
8b0899i5W8BLJG047ZHJuUYfGzvPaGa+BlCOMfSkJuXGtQJ7uasUPO79J84lpyR1l7QdV7+GTgel
bME+a65RhMDdLuZnH07ALLTCx1agrasT9wbvscWo0PQZu7ZjKHA+a5NvYc1/KfJ8jb+p8WerAZzl
ggJhzFODY7XDHXSDTap92qfbMd225fSfmIzz4ZTO9QWgRh5TJEOiG/Bab8tnlqjeOB27dR0aGixR
OpZxc407j6sFypkVm5w/0qtKGZ7GzyvoMuVAf03Ja2178A/UbCH/cNWY3ZK2NE0k5gbPYJheSi1v
b66rd9McQ3NILvWaEx+FbhGsPW66A5DA8lIEhmXT9fukIyKZBIsVp1Nlu6g55KkUpwGiilQqjw0T
7ACiY6iP+sF8bfxZaH1agiwwfq7b86AnIYI4oxt+3F54Z79kUGPrgtuMvu+k+PjXC7kB8DZP9kNl
+7alT/oasteJvl+vL3GSXwk0qcLlSmZPT+fyvnPCvh3/1SBoAURn5wgQ1N7CxzpRcqTFsPkLg+hJ
/RnSyZfouqcCoatd559ZGap5nKL5qtiT5COCHiFwwnhUmNKyzwETDgyljFTvIAPx6C4oDluIxSLS
oChkphEEhgcatuPUesMKgDEnxR/ymjTNgsODhbYkkM/oIBcSwSUrTwoCaCGXIm6x1cYWX81O161U
Hv8yP4XI9f14TnaiOoaN8xYi6TByy92xOB1SUdf8Yd6EQo+zbNGNmHWYCw7O2RSPRl8SroaHJK0h
Z26AHiOha3552DAK0JjPGbkTHqU70PcXuoxX2ubhIauTlv1z0hbb8+eU+AQuanHQzO7QXVt7MCwm
RgWVRc3UZC2Q5Qs1vSM6eGObuw/nMWBeMzfF4IrqH1efsrUVEJWA12UrqqkGbo12gHC1uSpxX4wh
jMpG6PkgbG0exleKG74KiAkSkQEoYHMQTddrlSbqFcxnh3dMif88hSzibxDYuSv1G9VSjA7TbQ9m
4N3GeAqCsBrb8wr/FSb29A27yKYlz03igcNemb23CGp0Z7ScsHpI/nsOps7ooVdeZHeyO9yCyNCe
mIwDB/19ipq5+oK8nJzxp+R0rHs1n85cfGahrfJELmQleHEhevGVFL0/XU3KTqdtSbbYqMqtWosD
AynZ/dmSrWmI+I6E2cehqto2cLej/DinAX/XEpyNJ0N5hQNq2hQ4r+wNj8YBzYGlRwmH73n+xpvw
PKabCxsMEBk4rZHQb2HTWwwfi9sBY9Ey1b5TCYf3NAS2H/P2LUsh4h5yMljmYPXGtPo72Zr8j2qc
taKy0+sntvTRyONa6aKjyQgtwSxDeuRhl6qCBeMQa4HzZPAfPVeMW2LPPcc1Mudj4XRoM/DJ8uBb
/4vXO6OmRAdNNopIL2C9rT1c2JLD2FTvo+NKgFeWoCLqHknXafH/OxtV/bjqJ3nEkOSxZwHQ3dXy
oeEeL4UZP+sDC/KBO0bYc2Hru0zexq54ndioi1K8nf6pxptMaoe01HE2Gcd3uqtMPW+8XsqQ89bW
ghpzn6yUQxunJAWT6G6WAq9ntqTae4zfltvkVaspMW5mWrvjEUCLKin1verdjrMvqWpTQY8T8cUN
17AWTW/siuBNIYpnrLHCFjP4X2x56gEBXbMYJWQ0lZd6y1nAMcRKWL3pdid3/TKUtaERm1uOijB6
oaI9MQo4a3LUAl6Sm2SjeKKEEyA2Vets3CkxTg5/PR9YjRvwo7fQGGoe3p3zReqwFiAYbEgbs+TE
hJirOYwtPkOpu78FxFayXJGFHtidlq4jIiQCRVxy5s+KlRDiML6sy4zrmh0s9CAFtfadxWIOybQ5
xL4TpTM/km3RNPKK42r4i/qNh5/Pg3U5o6Ss/vFaRLzRH/u1bmaC61nocE+kfswhz9MXfG/LKGfz
oGiFqBZv5eEH4nN41rTTL6Kq3XF3X6F4RB+hoXlMf4TmnGg6+QKIhxYBnuRPKJuqi2fq2/1+AvGh
EPl44gkmWd2eCI6DwVGpeO1FINlAYGftpG9HU/yq52vq6kbmrnLaBJ9XChp94dDMcHGf2i3JxKxv
CHdZWYUYG41Ru9/omiI7H9k12rvkZUBU0EA3GVJaMhpUPnq+5hAA4URKS7gcGz6G3+xBu/N8zRKu
eEx2ffBJ5nOSMgAv+Dkc8AwHNFe8rkYRyDL+5rwV0JEBlra3Hf9i/V74Q6Fyy75xTBzkJyC8UKR+
yiiLwnEEacLlgfVbgWfE25DOhpa8htXda+/fN8gL9pva4PTVQtZmoLo9/WtEyIdF4jq2mBzTzOiw
gH2hY+4lGX04P8mcKj1n
`protect end_protected
