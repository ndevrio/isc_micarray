// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Sun Sep 22 20:49:28 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NoX7amEqHSbQfye66n1An8Isi3Ik3hBEZgzWRBvQvrxKYmVDfXxA5rO6fnca+kUy
1XoeUHhAy3e8VCCS28GdwY519SLaiVtCym9XP6N7Co5Epgk9ZISULAm5CorlfHMv
x9o9zcjSxYuBt15jj8K1gkR10TpBSlF7LgEtN1pBdZQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13616)
IzUnM/bAJLS3r3tKZGPzHUGdDVogD+7+rExdfJKsukQHpZQpiwAR6KeyZlw3jg9y
xB22ZdtxvMlL6iyfvyBImY8n5ggg8w3OOL3eOEo2BplrroXi3aN0Fhh+Uoo+h3eQ
1ATE8cYGRiM7BC6gOFp/2YrmLnzr2r7SBevAwin0+jEUxrrYlIXOlV2TRVNfqbuu
/mrq0LSx9ZLBAaarUuJcCBqCMMYoX9W8HVOTzCyjN8FNuT1Y+QvRldPGMMvs4rpm
MwsbuowS2fDPO6wGIM8LYS1cc31MTbgTYpPvj90SZgBwc5nU2eX6KZgsrusdZQ/C
4oebUSILx78+zq0AdyrFT/g/8fQQs7oziCTKBBqBeCwEdSAFrMr7jI/VLQKVMJUZ
1vspVbpFnCWsYvMKlH+Y/S7uDq9C6Tmk+BX/WWf0gLf9IDX4Q2c/ls0ZAf02tR4t
zJy+X5iaDhrdLf5ymftiSchS0PUxRQCbY8AScuJAK31k/VOSYIp9v0qeFr5sZOLl
mzhaFJ+1NMD1AEp0R35/P4g1qMr9xqxBFgltqyAntCcCPQZQlIatrxEBD7bi9Mvo
7yVlIJ4sFF3RSlDrPAxs/y9gkT2fXdOpcD5u1TEpsQXuj13h4qAWMX5zoE/YIPPa
h5pn78JYFkPr37Ws8AQeCxyQmpbwTaiDng1zPOvxVMn+uf7xfuFBIwQDcwcQj7Vx
8HzyjNTz45GdN7eIACmogSr/zjqq3Itd2TalTk5I5nStXzz9E7GA9tOk55fq6R/N
g187BGapNpjTWb9PG8qyeHOiO9J+ZOz8qUGY4i/ffNsSlSejXNHP1t/5rTPVWoAR
XCaUvshqqdtdjz/lQzjC7xxpKZN4PkIK3edM/oMn1lL07Bi9BnpZcEkV3o97HFv+
2ut5sKFr/9I1KeD+dNQh3T05MLD39GfHeVePrk3rhKv/ju+nzDBU2xa+acq+a95Q
0MFRoyP9r13SnahF0GDVMwo+VKDumTrEmWYqneiZX/Z9OOxpM04a43jLlHbNO6o/
hf5hx55X7xs6AvNnYa0rTuoWg4/JMQRQMY5iHEGAtTq8R3reYeje6mMlJrYykrL5
+s73G4nijs3IG2ipflvEHs7/vn0ULiVr8scHpCm7IRl5IGfqjZDCToUntdZnvncC
mVqkGp+MC9TBdXSxNfI59iQZr8bJZUqDaQdHIRiSR0IGa/fmcNXx/CMTKCOi6U3o
TtbrrBJioj0brVg1UxClEePX0FlmqllEVKyaIN3KROIVj4S4wrta+jcssyro0kuF
vZRHvf98n/edPoiFF8uuYWNiOSSVioZ3cIb9sACgNzu3HttkAvgzW8A8SUGqPzp4
GVhRBeaM1WYrIZqrrHORVONi9ziBHVqZVgeGCd6e0p+E/686JRJDIS7hv/hGktrF
G7TD+OmDn9DJ6D72NDPxuoPqfVrb2SqdraUvk2pGLDiZ6I30a3dN2VF9GaSJTmC5
C2SklCtAAfoBrmmmZyIeiK5dUIeJxDJJ13Q922WeIn+lZo14mM2B7192aYqgPjAJ
fKvLb/GqHFArXUWlOz2Cw/Ga3VverZRSOR0hK8ZkdWip2ySmfnh63YKGIIyNZoST
jq4yWmJGNA5I4cNfs6CYkt323n520r3yjxn0G2iuFnUJ+rZjF+T7SezJH67yKyqO
RVKYIFQYQTkGyqtZH8e7Vd0ayD5XDnFz2vW1USyGWRjbjL1RnZ5T5tHAiygPE6se
pvBkPM9iq6u+QtwEli14Q0RDyp5MxqsDOq1jD68/SAZSjIRaJ9KS4mcUXhVcJU2R
he+J23HkJYBbn24tMfRQNe8Hkg/gm4Y8+bhQvAIPAFgxGwOZ00/LQe3b2tuohasg
IZvFeOJqR8khPZvgMZIDQGTILHMmDmYDyJc3sXPw879PrFJax9T/WnBd84fr6uXb
fcf6wofH30FHt8cdGKGaiXrWpNSQlYukd+dntjW7Y5+7uyGsm3kZZ+YBDGf3uXUN
S7/vaC7qgTja9dkbT36RpokaMxZ/OazXhfmGBOrbE5XgRTVI6FWgWs/Rx3vFTkO+
ATdpdrm1JoE3csssg92oWZfj52/FPtqEu4ZE5X6Q7WYneLsJcJaNumehSwFCqooI
HdxokWgWajiOgshSbgJ+t+lN93yrYZn7bTYHLIARukXr8dVNVXtehKClbLrqGZGE
p3YpBtaTJij2+EEhLmJxChvaXkxcTVzzLT14XKqAcBCj4BGzP2M3zNtf1K4N0upW
b70+NsyHoXeQthknyElUTCpd/BWJ/h9RfwJjS1Iw0Wk85TsyhDrWgnEFc8dJl8Vd
d87xJfk0jT2UMKdLboaL4m7FipArhfkRxiPNIu0UU938EVWrRaSadhyItge6CeUH
+UTa5jacCm+JSdB/ItVFsKE6gbHkODTQaE8+rdlTLGsmKIbWBTl9F55o9QoUMx9e
AmGiTB+gwGWjRCdwKBJGI6zfvwLTL5vMSV2tOYycfSR40MCUKeLqspBXnkK0uRMA
CSZ9ST+vFDpqojlpwVtkjK14YbrIUSucHqslXjt5P0ff5bBNP75rrCXFpB9VHUb2
vaSNepX9b0wWnklvJpENnIJy/OxQpl8/Wi+y7SvgQiTZYsViA1pxecnL2cWgDGTG
cUwnyMPx7OYGgFlStfHBGztyieWR8XYkeMzUTBlUcOOjzXV4I39oLNvip5wuU+OK
/N619hiofgDl4Zs1xKQTydY9q2uB7/IUa/YCD72TzxG23dXeEktGYQM1/yUzvEtZ
waQR7TVn7tjH+BrA0/Jy6v9RebL8Ij3aovZsu7bQcfzeSX6qyiSnzUcCr69c+Wox
kPL5LJgHxhzy2x3nS8x6XgKE8q/0qQChdUzx6MQXz/QGsTcxokE1zNwssO95XL0q
INMH0ySOopb/k1OkVfvNpTS07nXLyioHELcLs/Dggz5Bf1kW2KBjAu+jIKxrnr9L
gz6FAeJtSuOlXp465in1jE7aXyYAWwJ1vvimwR9AZ/hM1/zQ30dgaP7Zx0NWnP6B
/Ab8XtwZ6i5VKTAtHAuEINKSs7ED3a7GiiqgAF6ixjRcxRmhA1ACPm0TQ+TBsRiv
DO+DgjxaqqP8Hzq+j6/c16AWOidK6cfCWjQJm2l/6QxNXS2rDD+kh8djA0uMXVD9
6m+fDtRVG/AHs9XKiiKAEn7GDZ56w01L7YMZmCvMPzLM3ddDMcHkCwheG6d68H2S
Ke6M2NYjDZRz9En/aJZz3U+dIpxTE2FBb8KovyNV7JFqxR4sDttgyi6J7A1VAdWw
sIh1XnTjd+FQ2dHxeXJV8F4IYa7gOhAQSDWVl5pUvlym2ARQNlPxEPtM8bc6n4m+
OS402MrXse7vOLwAHXZfhUKnqBVRf8RzbqC2oqe49PsDdAIDHsydYBtkizvqSuSO
rM9Akc9kVnISv/ZSG0JWwb9hT4sgWAL0SSmzanhu1SGjm5Y4VR1VQ0DsjCmo31ES
psu++v0lTD1+GcDeDhgN28dN3SjWw8hqOYaKPKhp9w+QwfngT/wqz7Sb679vj86U
6A9JHHI+iyNPgeXIWG9HaxyDTsm7dsy0Vy7iIGQuTZppgLFSdw+qYO0wE0b2gIvB
eX5lAA13SZlvDPxl5GB6Z1aQ2nOrcxUDV4OGb8nsEgLVE0kPA54kh7OkmZEcX6RI
0Twk8c8WAw9VMBnpTTDar/1JMhocFpPN9S5GnRIWS2tlFv4YBwFFiQvdaeNhZYiG
Icoi2LOWq2OUn1MYxtOlSpYPe57RS8Ix6fIAKca+Kih9a6SKhDaS+s/NPsEvv1dq
MRufvpX5iYDM48GJDwJ78CuC+00UfBJBpO9KNyy1QFy+FrINzzUTZ94vcPl1ZVDk
M7jbyIA10wb5hwaYqPmiwAVCN6ao1TWrauK90BZXcC/01/L3+Y5ZIhUcd6ZcOlaB
UM7K3T2aR2+uJFeg0mH0rHB7y1KiufpGbr99Izj7vbdXZSKrP8wDCP8rYTxxreEL
BvR7ZguaD45A46snzHixEZPto7OzK3a2La/8twD4fJzGctZFbjEjV9VncTARddNT
xO/H5ySZzL7ZTp+vfIUuMR6bO5EINUPea6C/jJxNet/fKRQnP8BlYV5gu8F1jjfL
KO3cHkaVGz5fB9I7FTA9SdFUT4h4SRvKXWyOKUBj4z494zT/gEgebhodpjsXutGC
h+CadNimy9RN3DFQ5J8mX0tOaVIhSgy1huH1wMxgo8k5oremzZLotwm5xCXk0KsO
th7e/wS2sWEjW2KwCzzvTjEUQs2bifYcuNYaYad00CXBKNPpJw6P/KXzaguChNqt
UFmDLgMRqoiyaaaURd98tQCkrRBn393jmyNmjh5QdRPfaP/vG61uRgV1FbTHfhS/
jQsLRJ4h6jPZVId4JRleMW2DPdsJGvorbJ6lMEb4SDEzNALcyAkpSkeSpDaXviJZ
L0etiM4Wnj1hWN/Jo0CJ6BU9OdNwkUg9QQK1AHoEq03Aj95iCdDE8GxUtmGzqca8
t5Y82pjpfA4bJUDREqUVWf+DDPRkIuS9a1GJiJVP9phJSUESy9hWwpfH1TcSgMuk
SS9sLthNrUIONk8d+kA5biFGUeD5ci4RZ8wWgifRb9+3xGirfLsVgXXNbt/yWwMp
l8Ho4Jwd+oBlC9fJaW29hzSYCK9uyslMmY3tZmzefmnHmzBWgZKOWQ+XFzYLI3V4
urut9woenLekeNL9nWUGQvLAuDpP4z9gcU5E/ghRIM3Hx7vTyXXTMeRkerUNu2L8
Sozbl4NbCWLOWzprQkDKwqwZu60D0fKT291G1GxqSreosQrur0c+s+P3vrv8cNvi
mZUXU/WUVBYQTeq8yqTtfAxyiUwhXwtb4wGohYg4EVLWZ8pb6uBDCv+D6XD/dK9N
M4QX09st8PnbueiVCJy5a59x3rFZNXx5xUA5LsmZ9qo1zezth1E66REPOCpYzD5z
BxS1N6DpTzpCAXH1DHPKiv9jAYaue8l3jPho0ktbkTrrWux+bL4pdVUyZmTuVn4Y
2w2s49BgyHwNgeKG/i6a72sLQrohms41rDIovLnQtlqcXkh80Pd0MLVWUC9Uooh1
ap1uSR/ogidNHL7ah8oBu/iL5PC1W+dGMLbNfpJZnyOA7dnKWZcNhaHG1fjFLvrV
YhkqVndY99RYFgLmXg7UtWBDQwjawBLhv4qusxoAmqxPLa8M0boFSoCcORyVnwLp
geljGZPAfj1bsUeS07g4fPWTQc48JzQyYRGu1y11YxL7Cicta54qldofsTpNMmvc
3bdRNpgDLoUdM1KtwyVY8flrHO3k6EiFrQOlAF8lFvSqn7SofOrIsFmXU7lfbw1O
l+xG4Y2oj7lza2kRO5ZOdv3PCMb1YWHs6Fe5OVxVPotGttAy/E2iyN4WCNAc2NaW
T1WkoYCr0mR5YKsyA4pz9ANJIH9PWvcUOF/eMtMKYo3tQYkB8XsU4fZCSqz1Ok5q
vk5Rd44D9bJBLVIWcMWbVY5I3rOUIew0HbDHiBQMn4S62vYo0E5+Tu2+4InY7m/T
n2ml5+pGdZnK2IOm5VUibwXs6Bd7CRFS1WKsNawRCpeYRkPATzQbkM3JE8+fMfN5
zxGnU1ed4YH3XHlnlyX0Avzc8jHlsyXv9ZalKgr/kyrDV3nr/nbvP76uHBYLQRV7
cl+/92G1h5zepYSm47bSnTmzhPHcLFMvSNbnvVxVJlIdlSrs4iKSg1dt9S2ONj6I
N3jhfVHApvm4os089wuZRKmapKHqbu5t7w4xKwB+0i5NgTPbbnLmTeFNtBvgMiDi
cnfwL36BjLipTc6dv4s4XyOBhbwbZBkYrTJHmQv8Hh0gCHj9yUHjB3SXhDOUaw25
pk0A1Q8lkZ5roU4RPgBZOkbzcP9GADOaLhJGn5Xv92W0SKkQh7E/maqOV9CnKkV7
mBjH1K7geBivEW7LC03CO1jb39yErdiaDMy7IepJ5pl8BMN99MjmWuT/o0KAaynw
vrkkmNCXryvB+PQJalFunLPLYeRxHkksKZlJrqhrho1lu/ld852T9LHBbvm2vpKK
yzt7dn8K5VUA7Kg+l+p+3CkCPUVQDT2Df5nP9xVMycvdg+ko1HCvb2JJTVhHNqy0
CFU+gxYronw/9lE8G5biY9ajkRPteBK0FLgR6gT6HWedfJYSCA1D0nNYeRbS4V+U
6zcripzY+pkHH7KQPtMMBylNUT5jkiSTG31rqXbgLHMi5r04xsNg9tJ4Zg5ve2ml
Q30eSDAW9pYvVhQKWzFsBbtsgq0s3iw7Rr639dy/SEbbgRjG5NcfRxx0MTuFX0dG
yrbZ7PY7cKFHdG7ukY2/5fsGWKjGN+rh3li3AsRdi/XynvUUDLaeGEF+Nk00+CtD
E0v9e7EnttUPRN2jEdn1HdkyTGf/R7l+eTYFGgk3IwrE/EjeZqkz6r+ukihADjWp
erI/0Jo/Oj6xrlUEJN24lNjJqRQhHr8RWPbGMwNsgRhYOMa8DitgygHWY755JAJL
8PMaS0FIeDX9RtLzy14ANbA7gMuCizZe+5GTHVpwrcWV1/8ARC4uUymTB1luQDXl
kn1elDTeM6NvYhOc0zyvJ37Z/IIneq16RBHjarAEoTvKswGr/4LNVwUhT/mFPoDF
Un52VYj2mApql5k0Zjs8Pt0Fl6gbXtvAlqQcn1lmXomo6ESkEy6A0+c9tCvAcFYk
y5NBGZqrUlx0HJ284wS9hniQT6n+c4J1KQ0CUTqaXC6Cq/PuCP5G0KULf1buMXzw
Ax3+PUxTDhvuJa361R2JAkilIzMalMNj+KhhYbk6zia6KnZqZumhkzBGEZPUT1pN
EFbI/OpWoW1bMJU67ighq0EA4ULfE2/pt2egi3AtQ0s/HXWwgbTM6d2baLtLxjGZ
lVw3deYMOiBOa78nfodE/CiBZM6dd1l14H95ulvMNLnyc55ccOb/uIgjgaO3yT9I
5HHpCCdpeMi5z+HFwPSawL24HLYwXqlXE177EQdFoSX+ODs17vvUyYbKu7MiUbM1
1h7cxQOhuc4WlxjikTxtXwdp9fbC85K3CmZpeY1DzAbN/8itHNvRDADdlav0kJj0
iuQ9sR98uFcdSZiqiA/xUdQt5+77ZDRzRBHn/8QLyf2blMsJReQQPkQlns1ote+T
YhjpXRfnFWMz2g2xS2xM68aAJHXG5xt5jORqI1S4/u7RefSoWIEy7yS/RiB+p6fa
QlH0uL4dMs3z4GZ7TP/TzdAkTmOhheDug/VaLswalKFznzuA6eOvYa4j1M2rx1gu
dLdhtHSGWNrs5bcv2bgycItHDzMy+fICUekKqAIw4ebLkpwrqTW2z7TtLSLgoK1F
erS3RQKf5HLuWyQHLKcRCYAH35fqKBC7jb/ket0+aEF+xIP2/NW+/hTlGuOVu7Tn
sN7S6Y68eShtXVf1EStORB2OD9k3T26j8qyS+dHqW+c8lqcVOczwoY1nPhN1f5zp
488vHSKf/ik8EoOPc1CCH13zp9EMeFsNr8MuHlQlX+HfJKyVJtyixEs5CGMGFttk
Hsap4W2CJy43wjC5+6Z+ydE9eLae7G6HimWpiv15Ie/0OlWtYrKdLSDgIn817QLy
lJBQQDc0FBj/fGAXVnlfgTEuYDj5WjlpQ7qQ3iJDcI4tylmcdQT8wM1m8O1l/3fi
J3jB8sp4KNzYlf7wuncr5hrARlihO83gowdHNBomlC9XzU+RJrhDsrOArVTwQN9R
iiFRtXm78PwZJfwOTmjMVoqglUq9fpGIX5GYKhlO2t8um55CTuUkgsBrFDUZByqT
PHhFK9ntn/oZrOuE0CMEd4Xisewwyc+lYPhPYedMhx+VPRs5+CBu/ui88ltvlEbn
jCz0EJ4M7/xVXMw371xgzFP5f+yRmFBbhzthpf15bb5hxz9GuyxmYO9eKxIW0aJ1
VitriIEa6J9yzp+UcxItA/btLV0YUzDEsbNjV9WoUA63UACejUbYkPPrnLPJYxR/
5qDptn+bz+TXvdOfOWoRpzQNljzy38vdc/QzXKhIxgP1lt8LxIA8+bXapMxQ/6ju
E4zYHTHX4F56rPrB4WdDNI2YQvYk0U+IXCWfkVOwlnI0+fK3mxV1Mpze63/I7DBV
tKsYZRAXobyd/Po86Z0abzhvEy+tqeCa1JgCtEJ/7Fq9+QOYp+6rnGh6QZ6q+lV2
eGCgJ4XdreYkZeZ/TyfseIkIphcwJ/YLFUE/GgAM5mZjhOgk5hA5YpLQVBp97slB
SBEX5WgFdWgZ3mOT4CImhNE/h2SVv4kt/4djG7nJDjNEPcLjCgW48kNk5v5CDFIL
hY42ucbQkZ3m6u5Paa1qPwXlurlH1f3t8IQsd1ndnPVbyi6a6tsa1CIp+8AB9S7B
+8Tq9NNWvjk0Q4PUe4bj+MXhT4UrxALJQJ54xraOX4IclxKf3lTElSy0sIJo9ypW
DNek0bKYOuy5ZiuHPRBKOHhKvHvUQIZ47KktGQQHP4qY6CFYYdvaC+vpIZBpDnwK
lKw/8H8HXho9iN9014ZcZnK2yY/QwTIWcAuRJAHZ+jZkcGs3IjyQTJ9Nrd4qht+x
KwmawOJn3gntxS+LZIDHGdFZFXNng+JayaUjhZjzc7ptJgV4Izds2XU+5OD5eXwp
g+RRWQjMnD55Duh4pJHfqpcr+BW1aA723OsgeIae/8sxIlSB23GPBTTf9hlld/ut
MSMTWvRmOLrxpF29FCmSGgDZ6D6rofd5nKeQvoEKXaWMDWYYXI11JDq/HkJqXx6t
hL0gjiV6GM7dfo/8+KTZUMwT5oFtiMDdNSJB/ZC5dJ2odGJMqqI+KyMPA4py3ISE
z9B66LNOCaq4pLF/i4h3XC+3kDcgn6mpBQbHe5z5ayDm/SU5sF3aErPHfhGUAJeP
0oDxok0224YKbA6/0s1/Q7zBHxZyQ8llFw5AZTRWQgYxIIQdZJpCQIhjkPwqSRXX
gkw4tXkZOH6/hb1JRFrIyHN/TKF2d4WwtQJH05Vq/7j7G5RaEhueQOHrK/3ZcrCG
9w236pfLxAsFEOWDU6GFd8j03v9jcp9iTnazGUg8a8i+7F9YgffBj6/nF/5u0U+I
t1+G5/4zsihv5g5L7eH9kzF+snd1Y9VkfBx8QooQDdUOkcuUc+P7cweSmCeNPsyG
bOwI6Iqg4MytU93LtQ+5zJr7O6vhpzA+DCDiqh8CFia3M941wpWGC+RZF0W/KMkd
Mpe82ul08U143BNlsz6y9T/JfFej/htMNtGS6m+P4k6qw0wf2bj19AX9wfJD/4oZ
6DGHkM1qrcoiN5zZQCmu317shQ9LLL/erQFHJCT+sz4hjbMoPIC/m3m59510PqTT
0EvbE7ol2qXdVBUihgARMOZ6k9lHdq1CyMe/Ot4Wx4OiMmXiplae8f4fz4nJZPxL
gUnKFkF55K+lpqzZej2NBuVpEQx2LDk1LPTdpSvVkazAYQ+y+jR8ODDBNV4ZmkTQ
jWxK2284MOCjo3zks6kwuQnbF5vcCNXT+AucoqX2bPCyzbiGa+HTVKUX17ImTheg
ouBqzlLzqxC7GB7AdQn7Djvq/lzpsVT/iWHUI5cqoj7OLBbxt1K2eTgmLcTbsW+6
abes73UAL7Y/7cqOcEnSqUGVAhS+QKGkJIxNUlPU7xh0uO1s4vXI+fxKn0XEOAeR
eTq2a+B4+5S2loscfkUPnd341CNp6qa5Opu1/uxUy6KIireKuNQmPodnO3sGOe80
EfyYeEbfw72Yvln6FnKp+PQlWaPsY3Ia6CYtKzW+v1EQ1Rl5U+vnmqrczb/t1N3s
65RQSW9oObLufc9BDhw7L5olPdU4IvuImetZc8SBIf0zCWSsnewzmn1RYVOvYvBu
0Ik1DJpEmVY/HWnEvS3tnGIsRPSmkhmOjd+VHETKcBTnF8speSkbD7CbtImWUyj9
eTNsJHMFLOyVQ/B/prR5OYvXG8yPMQ9czvtRjxf3OIxN2JvQpDZ3t3KJBV8YSIha
ZlZvgHw+QEE4dpr3TEqyFLpoU2SbcfbpYJw1Lq6IHdXeVfhOPUVg5qFrBglUIPYN
NdI9OaWzSPLv5uccVZE4KulpN5mO4YalDxvvDnFjYGywWgr9yKC5gkDdAN2zkjPP
37NLsKy/EArkDPcQTxe0LPN8IFjUhbFjQ7tPuvVVWxXkl93HMyrGjWrDSDUXTEis
TpMv0XA+thl27miwC8xS+9qKWgPpOTmf9DfczsLguxBT32AFHbA+l5La1PP9iq2t
FPI2Gu1MX2Xf8ZCwUD91CtbsqzFwtro6fEIRUyNLupeI5n92m2glpI610T1a1n3J
Lsr2O/OSWFpgHzBO2UIIWDNG/1Gjg1UcWjnc5AutyxaxLo6+9ZNkgldvRIFZj3z7
ZLiddjDmDQCGoCSgCYb3bcdbyKdcRU0+0BwEkkabLaL+9lcYA/2fecddAoNBHHXK
HwSEg10pkx9I5l/pgV4+qrHczH6TH6Kw0+w9ATmlH2XhMrVrzDuHJWGv2ynvr6AX
K0EzNi6gXu+vfDDygbXRrB8b4Ydvn1BYUyyhtoPybpsxvXLoqycgcahEo8UQQWQc
wzhoR7uWE3cRc1qiKE0Tzy6yyJvd4iZCkYhsexnnJPwqwfbKi/pLracHC/PM/Jny
B8g0hkg4VUJVLaarC2ib/xpdDkx1JTu4YUZ8vDz+qfMU/7/5LrJ+sk6FYrChStlv
RM+SYqKfZdoFBV7N0tyJRkRrXSx4E0YGwaPDOsKors9U13MoXT1qKB7OV+eUQthP
LLCla2/O+QkSpsfc+GtdsSuNUQ0s6rqgSt0iv7sSwdceHaPdEEV+C5jTS5HHvv/h
SiLSSp817TzadFc+kE8PEoi2+ZiJ22k/x/sGC0Q+VayuYZbSlzb4pzngIoyWR+5M
vSsxYAsSiyoCi5jeKB1vxoxypt8cWPNT8nF0/zaPqBXJFerN6IDWLbjbfZNzAGMe
kV3qFapokNihimPTIRlr5QLv5QWKgP4kaeRF1NtahEi1aO4DT824YRSCmiDiLUyG
ZpawJcbfn9ZnFck56mM6lG4oXgqKg3YeT+6X09fPd/t53Q8FR0Uhnwt9EjLmKQ18
aSkkzahje9CYEc2V9xDGoFQROai/bO2pZ6s5nMtY0pw3jXrEH/JXlqpIGaLLqzkI
i/Eh+OofkNZ2AdrADvaGxnoLQ0rSo6fS7sP4fjRS0cUuQrF7TeAKPNthdIdpz0wz
HoQgz26loYJTDQLnW4LVUdjVUHtpC1FEnabg5He7AsP2CYjUbWGAANwdBJy2YV5T
SqQf7J7ogNgVeZvShN9ntdlO0FeibHRaNIZeEkpdb6T2Tp5oDBC4i0GiVSutrJrQ
xWLwz3mX0L3bSRuhvbNTFzvrATtRtIOg2qTQ8itflUlSCYA/TA6x2D+iJ8mUmMxo
ywrGv3qa5EAy2RN4cP/hJQpEYHT5IWH24ldR/n25A/0cz4wNoNAA7vn3QQZ5W0ZM
moofAej5ouChsrdc+bqR9npVxtCUQTo1ECFdlCWb6fVvnajshoWcwj7vpyGVJUY+
lVF2SBuj55BYz2NyMf6e+w/JHeNeZevs5ugTflDzyTvsQpd/sQNoFtFEiIws/YIX
SePzOoVOmxyR70xSeMGDkoEPPMxaQ+LmysK7jKcmsuD4oBDQIyoDbjon8yh6GFVg
69u6D/oQ7wSjIYVIOODUda2EOVs8zkgVjGAtDQy6VsJDOP1vRrhDWg20pSCtolYv
taB0N85/1Re0nEVcrRwM09wUpw+7DHGcqZzFvWkX92rCh57dBR5g/qVkUoCJrIgG
PAeofkkjWiD8U44esUA1nDnl5FvGri0VqmxU+CbeEJ8QOyMv2tAyUmm/wJBtKuZy
yAIYIVuXe6NTgux+aAhT2KhUufvZNE5yZm+YU9WNf3iWp3Qn1w02q753hFRhLbDl
SF8No1NSifE1jNfJklyMWNKW4s4+0F0cf7oKu2EopgE2m4rJiRVnrjk7a6wgzEHf
dDPIdCmshJrXBR/Fc6R7YmJBFVUGoX1wyYFXQCPB8tcVyiFLhVQ6/Gmq9zyLAhyM
WnDHQCkwdg1aUBiZg6x4WseB0casx4n0U+10KVtR3bsmFcd4CrB3xHWKrimXGsS+
KZ/oy6y1RH6djDquJdWdMB/JWibslNptffGEAYPYujCiZjtV7miEihh9RkBHm5e4
LctXgko/umlXOIdY9ucJj4ydp8yDGdayNXpIrtceax43weZM7eGZRlC56IYPm+GC
EI1aKYBHS65/8d0zXTmvEvdslfA+gJyN6mBb0YNVngtwAeQkc6iLG2tvmUzcNV6m
hE/o9RDip9ZGboOaXgOHJ6/0FMlzv/mlqYUSjKZIWev9/2HFLPlAxpOd3UaJKLXo
hTRR0MrPd+h8nct07teTbVknJm0lUm76KAZW5nhmXEnWdJsnH7IQkKkEWlCJUbiX
AISxMt+bknyzb+wLyhddxhi/wA5sP2531xqlkp0WAGDoCzgxqa1ZeKgfNb2rYYWf
hidhtOAcz4Z+L72otWPIrYoB7LoHnzOxS1AoU1+4GC0DcJqjkpSn8puZ4NHChnHp
o3o8eBsxESnFT6Hvl66KbNH9CXJQjlKZVQJaMSCVTkGoUqxXIuSE1wc1GZyMWaNi
zJd5gYKJ9VXuY/ScArjEsmIrKSJOi/48G68MU3uFGvpi38A9Dk7UXbrkVaAla6wJ
EbCsGCmSUF3iqdPhM2UdPGRZ2jmSULGu6JrE/6BJY1zMUzO/cd7xO6NQ/cw5YUJb
nIskh2cX+T01skyyaMHQ4cvCMb5CJ8Sfu4Tpm77o45pnSiq7YuyswsX8JMpTrnRv
hRJuAFJLVtrMYADjAgxbfDLqlYnIUSJQ5nommcwXot/XLDNNKRw0TZ73HE8zAOO+
41p0GKioKTNgH3exOIRAJm2yugJaMAYFg0scXTOa00Kr8rIny5y3FvDtDdjv5gdh
0oG0JvyoinlHqi+wyu4sd/zH2kjN/vyjfwaoUPXPCAktdnehfLGrfdyrQw7lgqQV
onKIfPwwkqElhLkATK0lzOYylRCcfkulYSZUQfnQdGh/G00Ql0B7ooonCF56d2sT
0JNZ9HdzjlaMTm/kY2kK4//5aoDp1H72wR/O+dpEJcg6F2ZMRY7DccG0WZ0VCXvr
otOZfgt/DzMssMCTy2Jw0gj2gUzCUb2EnANJMpl/EDfqs1pj5B4UfL4DIFf0mg+B
1qFYoi96vSdJsPuwDGNat+KbnoaE1KNtKHND0v7fRlj0iRb13RMVsXz0xZcKKJ90
+899A0RQd8zD1AJRf6ND606Ga5ZRkv+AOEmGjEaqCa2xMqzBRBFmnDcAgGfUeQqe
QriW/WXw2mH3bqW/q7b6+Guh6jAzq14i07Cqb3zNADZr7qvnmtVwwQn8C1fbvx31
A2dgbP7zi1oBV1o7QBOZa4zuUUV53EmvQEVMcpCYZFLZbi+cyYaRRsmDY6nWGhMR
rCSEGWqHa5bO9HAfm+35yblZkXOHIBxPtQDWvN80heyFXYX5DYiIS6+RIsmBtz+r
PkCA5c/4RPRBHvlbvx/gi54LMAGynVqxdH6C/69NEgZ8Nwpt9z95y3dTyWbOQuwg
/4Li3h8xbeYvkwBNcvFs/w5rvPwwQt5WbXN4+7bCHiIU9pfDZXBgFrNMgLAHCPDT
/WZMHa1f/qlugX685KvC+e085RmeqHkcVt/QrbTwCXZNVsE7BnaLcoCqiBBbhAyc
AfA9eMAerr2aVV8/zJmjg9nNTXlbaA6jz6DvZk3lPzGtOVjpV1nhi7AKEVDyOLKi
LZQo1+8a9Qc4HrOkXW43BupBhdykM43qyK5yijfuHoLBwKBJ6tspbaoDIJAwCKmZ
fOeWsH1NnMdk/Iu7BXbwUSO4FOtMUK1TXaHj/Zi2B88Dp4HIWUD9951Myug5HGhR
4gM/NQ/bCK+zRyBTgWJyzy4iBF2zUZiq8RRV/vxobXgVQ78sOJXnSwkFKeTxkSOQ
PpZZ6xUAQHvUZj7T3eHUrJ8xF10FfLljcN/+7ezRKmXD9PUgRqYNaVb23T/+aIQo
cd+25GxOz6AaGFrVQZyYrwf32iTojSMp+bwZeK47otX2uGNN9oO/Qaq8AKNmOgir
O1HSF6pYlpRz9vUOjnhbivepQMy+xbZzYIAQpPNtdBMMPVRLzh9jqgrMsE39Iv/U
8VThk2TOrS3aMn5Rgezi9yWB8LJdLbyVTTYA1/Ru0BoTtAajXdY6CJj275aYTCFN
NznqFYQCwyq8az04jgTYkQS6jNVteYlTjIa8EhKHu4EYV+YLQB5ZGGyqk+axlOvt
dcjriQhDdgy1K6yS1IologB8+ZAtogcu2GIBgH3N+v6I0lw3N+ZVKcgVLrqi7rJl
DM1KEwtAAh+u263glCEKJsCupW8m59zCSQ43vtJBV0XT4I6Fer9yrRxlvqrDQWOx
W2RuoPp6y7Aky/JGqgeVOg4wS+koY4SFJUsqAYmrYugZbkPG623elebx403HPKbm
zf7dRh3TPY3t8ynZkc64RA4GVsgw9ybNwWIWF/4ZXZ3om/kNWsEJr2DpYNw1yX+t
ecdYAtqmVd6Q/OBFAA2X4oZoStwz3DeOSDGfeP4e3EWY9dfGP0dk6OwMw/vmFfWy
SkmDFWik901eeZK7gWDZsC+N3aeQ/cUHmVjiz499cE4/IdFpDQqS+mxNUDSJyoDE
Fm0UOcp9QhUEEPRgHKJiNVbLKesj6ODQ5fhnoKxOYoH1//yIw+rYz3w/QG61MrNb
Hs91Rj6QbFCrQ6U/KRC2RRwUTSyaCYPDpoEg25hptoDLHiPrFH7o1KTLm5ZIF6Gk
Fp9wrqD5Owms4jbYd0XkoMw8KV+rCEnrXmm7IbW56uBOCdMXpBAnr5vDtNmhHhxr
o+ZeqEIjReUd3Hr4oNrasa2tNBKLfo7GobBrWAGTYmi/ztj7Aj/odamotFYNHcgI
NM9hBpJtF0MBFoQl9RB4O+wtXdXkh2GhYHcCeHSn1TQFFogJO3Zi8PHoEo96nkIY
8QLzNvDKY4qpTfqOyPfibv5nJzkiiMriRxZzGzR8f2aM7eRdAEnM25CbT/eGu9nf
D7FJSon5g9H/cjP6RbzxFIXAs3kPpBJfLNtKz5k0GMn8+3UralOoKCAcDwNebH/Q
AonIxw0oPGTu4ydH6BMWEf1MeXYOSZQbhSUiDKU8tF425b350drl3nPalHGevyPm
9ghOcC9cRmGY6slltTYS7g2NN/iJIrxV26rOBFFebwj6RwQf6euyn8z3/IwRgxIa
VSsEcNd6HE2J984r8V6DZUuUmRbLJ4DY3seS/+IudcoguaBFesdO6XTE2Q+nI6Rl
apByYLFIz4BC6SGzmxMbRlVN3cnCKtFgBUfqbHDwvl9Vz2QoOtof33deXOgpa5a8
Aw7mHDpIiRZpRAaqZhVvRDC30VbNwlgYKFkZhPcczXIaxM6+62RGlM9gNfodcZSf
xiqaUCdKX21I9lZeg5wypM+QlMQcpq8sSzCmZhy4wHlzMuNGMrS5Vx3VmrN288JZ
izaODzf5MeyT9H+ugq4jHjIQQ8fK6bQuBGirmzomfR2Y1zwp+3w3hQhICKcCmHM1
F6UwnNP+RfDLw2rIIdqKqtMINKYJCpegqGkQQVlCtd9nYpRboAIP4rppyLB9CR69
aVU1jSFxX/zSObNy+0lrdfLGLktwLFixfC2VnF9VGEDIrp26OBf54u8XeUvqK4xY
XtvWFF0RCxeP60miXgYZoFva3lAzEO/G/yg+0sc1g0+WULl14nPZ4Po2y1Chso3m
C7v2UrdOxYmRQPm2AwS3hnEl7e/02KmDsc1GiMbTK+7pG5RCAVc3oGZ5lsrVupK1
kqjvSvJrdFH5zpQYZZo/SmsLiYFbcK9qr90BZiWi5AjkqXE797hPMVgu5VR8y+PB
flrFnK+Q2SQtSFa6HkP2k2ccXEJBaqeIr19lbEsxXPhG94DGrOZ6sU2xvAo+4Qjy
BY3EzXyrpXUZdk6l9KMOIhgd5z7adPEcF2w7lq/nf7XcgBbRsptflyT79S+xWraD
8oDBDb9xyYBChLyaAKxexGr3dY62zqGckxdE/7pBlNj25GASLwKklaBkupO17QjZ
PeMtofWnLOnLvIetvogMXLyOgvDfuP5lgn3nVyL+gzlS5VYyodHaQ2tht6yBgiV+
9zcZoHEf1+7kpDfQKMMKIvcC7Bbd1noQiANmDlCZuJdSpJoBeg3tYgGzqjhNUDs2
cX65aBJp1RLwRo7i69dYx9xzrxJIu6sd1XoUPrergmjBnh/v+eX1qxbdJznkPHWf
AqdRu3VH+W5aI2WwjG/U+IIO+wbFu2womNlYb/SQPf0LPZOWwZdBa37D+R/UYCLD
y4LMyIQ3zKpp4x50rRz9uXYnyVJBaLyLmQB/NkXZGI5K6px5A4EtX2oOy9U6Dv//
9VcqZpqaQ7WvLDH64TNGb0UIZINEjl+MYTRzHeM8g87cJBDZihF8z7dj1qO+OhkB
RZXIc8sGyniLyzkxDFCtstY26/Lg+/6vbmhmCtLUYHDeXfNFJ7lWHs5jeW5HcwZ2
3/2zu+Qb8Ec31W7hU6ygmMrGk8gDdbOqN+uq1KZw/6AzZp6Te20VBPz5LsMLDPGn
DDZnINNBHOa7XpEbUqgMMCJ06rc/vyZurnuCPp6QSgxV53Ns9V8KboHiMBlOy0NP
iy9dbotZEi95aNZSh/Eg0tWO5pcHhaQfqw8t7W+d/uRC9m+K1EYVlojLt6TaKIlw
SltG7G1i5lHoiVy+RyATXIHNMYR8t4c6PyITGjh6YjJ1KEVl201CZ2PHo3Wq5H8x
m8/ncU/uitTvEVMAf6j3Dyv+nwSHkxlHsv5QL2A5xY7pAOh5yo4MCSEiMPKCE89r
v72JuvYTrhHtODrYbTVNqGBP5tR0fwr8OShyI4lCOban/C4foAxY2BCdrmXOfijG
abtOCOGdmwy7p5Ig+g76lR3czhYTJ12gAuJzRc1UWNCBw4rNySa+5ecAz5HTcVWx
EGhOnUCa2wTr1j9F+s3w+GOyOumNCCkwsLHXDsx5CeJjhiMPS/WiCFo32NDOkR+M
4G+5Jv28W0oUzpdWX2FK4Mdfk4no9zzDlMf4li8BMzg3nnTE0z+Qs/pLVMixHovo
mEPv7k505VyQFYlUcVi7LRANjQU9FXeK7ktQ72l9tJqgYAFoxn0KUYEczt+HzxOn
j0cWbdgyHewm/WlEEMzELdJPP1xWusTyzlmgBrLqi5OYPLGf7jOp+o7apYTaQzls
UN5DHfbwNBdhfrA0FXheInWu8+PGJ0Z2kXoKahFDXE0VurCmrKL9a6nZQvDV/1GH
TtjXthejzQcggcle0A8KUjO+Oyz382TyUHDHhUUR+XZZiigkCm82tliDwNhm/4hx
NKF36VcYISJU8vDSfQXP/9huqf8wNWt9lKjp/XLmGzE6Zw3jdL/tz2lsmx4djw89
b9boezvq0FGmX1DmlunZ9oJILLcl4SJe5l4YlUjlIAUG5fKPJqp1uaArAgWHgBy9
4B2Mc34dikHLMYXoNK9WfyL6ub4nC0kLVD0VouU9u1kIpgBeTxFUEdtAPe6imek5
ipT8nQR0Ws0LLJQMlIsefBmocfQU5+k6wpLnFVACHN2TzBCLs+R2d8v2y4YQDWO4
22fmzPOtunl9189KA3J+FfUOYBoH4icTVa3EVBq3lrJ4kkqrMpsm+u+GvocL7gPz
HzAgfnPDRFya7x6smiw12DVneHSGRmFLHAZXANpNNUaQTF5C/swakhauwZKXrLlB
BMPgDYu+wzPTDXAIDG2R3aKQt0H1Tk0ppCKWWH6yspuVAeG4zuTqv6PS5JGneU8R
bmC8VzH6ScjVm/iQ2HK+i2tL/Y+q9l5vgPSCi9mSmGfehCoSw/D13uZXJ+wtgpbK
+4SyrMmeaJjYSYIoFGjYn8/id7NWEqISv+/HXtIHNNULvZcbFfWJrR6jRAcsYZGd
9/0Xpa9/Yl6t/+WSY+tqu4xBZDb/KNwE9OyTbd1KJaNf+S6zG67kYSUng8Y5Mu6B
JAWZgrygUEFwGPWNk1pOLRiHFCTMpjuveS08mtM8sKPFbaDcnxj93C2mJN82vuIa
JRrgMjkm9rLM0uOvqZcJlvaBqRJLBSZvm9qhM43311g8PshugIPu+ce3h82/lDM7
t2dXWagnHT8nfmcgd2p1kZj0/svbYOt/j/lv7rpdt+qMNYNQLG2Md2CPXrZCPN8y
JPb/3QEGaHmBxNXskWlT0F0fuvm+H/wpO3MehMxCOFg=
`pragma protect end_protected
