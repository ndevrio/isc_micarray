// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H)5'$OR2D?P'G8TC\/EXTT[!B0G;X>2.M'S1#Z%SS[O80!;!1/F?KU0  
H_/ 0V4>TWV/YXZM"8)Z?W0)-.OEY>1A3][J3(BST@70>Y7:8=:8_80  
H<US<1+ "3N8]CU(..?Q&8)?=_$8!+[IR7%*E\H0@PD?IMV2I)X1-9   
HM2)8;FJ" EL@*9DV0,)X>8)#_>YRP@17LA<#L[-QD7GFZ5 @X*FJR@  
HI-P)UWXP'B)#CMKVN(*]@1M0Y6J/>T]VB$DS1\HBAGBT3'.M7R-$H0  
`pragma protect encoding=(enctype="uuencode",bytes=1264        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@]N#OSLL7>/0Y2D\4L/]'/]1&<:K>-MA65QT1@E]9=WD 
@-E)Z_<OI[/2@:=NKH/BV#RE$QC!<F^@]0R?!>BZ82\P 
@.'+FF^=)X; #)T&\P:E4$\*ZM$*\O>L9Z)"'Y$T=ETL 
@'2I &=[AQ=H,[HL*J#QEX#<?A0%[W?%<^=2#F+4SB2  
@(]'X?H'XC)####ZZN-%^B\9Z."(PL8UGV-N8=;U-RE  
@VG)V"G :$FV;^TUA0T+ITG2AJ.^07,%M<9,_ZO-=(W@ 
@.5?[OV;:XS(]"3;TD*JO"L![APVU<>>Z-EG2=Z)>-5X 
@P7IH33X:?%^H^E/;+/$GO>B'&EQCR(WG/2J+B8LZ?OD 
@E#4A@%$J43W2@XCWS=MNE3%3+^:S3]62&6,IFF>5&(P 
@UK+05=V%8T5"B85><E]=0Q:.UOST3B-DEL!K& ,F=R$ 
@4VB$KV$(F%%T,PP07X%M0(M-=S5 W7XN>Y4+=M&!L6P 
@C?#K!C-^82\PLQ5$0E0J.#'VU8>Z94[%.8*(V0A#7I8 
@W6)_;8U@5UG\LW0EHEHX5'S@%2^&TR<>B7-:201.>1  
@$63)Y7<=E]OMYU,=,)0W(Q$;&Q9D&,'O_E@P!NNN*5X 
@'LU[XTJI7FY7%]=-.U'&GO_-;^U&+A*+*/2U_59!ZZD 
@R4Q'DK 36%/W9;JBG?*AXOT@8BYS"JJO)8!_*OKU:S$ 
@&@PZ'H#N] =N2>A(,AB*B87X,9PQFQ"2(I5O1D?R^,, 
@3^_^5)Z#\?=Y-E+I+R\7E,A^JVDJ9]B8 V>$U;R"@&X 
@G2_2>*!"#3 F]+JVZ<!.FO=I<ZAEK\,L<%F#"]Q]]B@ 
@PM$D0]U?2IL<N[!HU^ Z2@8.,GDWKG]/:_P*(;M^N4@ 
@7'7S6D1>JA+.]S#P(K(F)L?^!/W;":6=#RJ-0OKQS/X 
@;HLG\MJM.X*M_F^!*O?\PZ'NXM\4U1IS:I'-*9^VEL$ 
@$H5,V'G2F7X%//91*O,]*]=Z^'H*O8(/^JTY%W9D'?X 
@T373.MCY[CWG#5 @KY#  SCC-+$F0\-KL>2[6P8B'1$ 
@63L7!.<$&8UPM6R]0.HD;$, 0%HB1C@70^@+0V'(L+( 
@Z%1!OGOL9+DM<D=+/5ROUK3:+X!'-!.X5=C1>U)%NYH 
@Q R&)VG&!BNMS6N:;IA&AH;[LEL'D<^L )[R"BB:T\\ 
@D'YX)AUX,$H[_RD]=_Z-LK9)S2;WA>[(F<^"W1O\]70 
@9/PU#K@LCD-R<8B#'HRB_9$8JWHE?SX,ZZ6,7F*W7 X 
@K+&N'&@O9W=G]Q[\A>6]&QEL^;S T6L-&YTQ/HKC',8 
@T&:%?@8!(3_Q#!=%#^]*8&KO!Y2DW^:%A.F7:H_W#&, 
@NA'<TW4ERXT99C>'"3#R]?M$/8_AGK_*=?%@+;+MT L 
@H  %Y/.L6J95LA,@.[K=:]TID-14H\)C[>*_3T19Y_X 
@..@SYL7Z?/2/CFL1R5-S/DXT"9N64DMLT-^I!4G?SK@ 
@UGEWQU,1;<L.9K>J\<%&=4K+C62O+\<K&/3D',"X7U< 
@V5X63(W(^RD?)$5P;?0G&LS_<?DX;(^9='/)9M0>\GL 
@]0*'3XYIYY3B%-L]X=.'3,D$KFU=%].RNO^%5^D_CKH 
@<\O,;AN/X]\;ZU04C.,**AIM*V,);(3>"I>)]ZQXD2L 
@#=.V9GZ5686>Y0,ECLVP=]4S4D2F/W=)7V,G6>WKX,< 
0S4BBYR_?+DV!5AY:6])XD@  
`pragma protect end_protected
