-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
dxIBQmRhEJ6PpGMzhKLMTdHlR3nbtbx6Txv5bOhhcrsJPbkYYtblJRS5entPuceU01TB1wUcvOt1
ktUjd7E6IwfYbTRaSK1hxi7E0bsboyG4e73FGDvPcy7Trt7SRECkRjHPiSWGNXsHEEEIx+mwQjFA
dsTRYpoehkKa0+je7F9JxiCVWm4ijTM6YTwIQJ8FhO3UedIsuW3JYMWnh0IudVpUYmMJwUmlPmwF
WMXfvqK0vOCF3LT4292jbeLhoMv3dyInKY0UWv83e0BvaLbP91oTdXo5wjoVurra4uINk1+hHH48
s+ALp0IllI0hFJYWdBtxRthoI10fzOxBxy7BRQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6496)
`protect data_block
pCgFCDQBPDRBqVpQwaz3DxTgwToo9I0HWgh5CLz+JPwA/3MQDZVxk58TSSovx4KVe2iviVJTU4Hb
3xhr7cUtS0mFTWda5mml8i+BRU0bynO9ylqFNyqqPKmW6DXCOQBoDr/4zeVPqIq8+XNnnXVDcUL7
8HKtvzyYWBX7Toe1kRYlBsqul/mNAnfBlELDUnvd6zc4BVYPClrqeIntqAYwLH9dKx+Sbu7zJSsq
Osqzisvx/oju082jv4tbAzMGNfF91C4aq9qoYPlso2ZnFscmPy4YGxlSEQzUwraeGOpWyJYh2X/r
K6Aqndg2i3I7vu+cTG5rWEXD4XTs0feeGgV+imZ/ICy9Lt+DwzFLddF1nk6mpPcJF572u1Xp2nPs
gEIZaWcK+vJP8FWFtbP86dM3hjYMax9l25AiW/RDpAKtc3aerEtFANooQ4A9bb08sr7B5pdHwfkr
uMHbc3aN3WYEXr/Be+tIyc/8rICK9Aq0jXggrvcGyeoQMvvQm/XpPrhp6TnUqERcr95dnghdCqsU
IiHpf6d9CxsEqxmtRlQH84RJk5SQpu2M1A3KhrZIhiql41U8U1Oh2Enzy4/lRW3yP7TOdaTcX04P
uACUKnh75XdFLP2uVsvAfFhGwtsHSABHXJlU4+xS87zIkfgc/OBy6eAZ/06/UtOVrhK5giYJdxiv
u9rRrV4Lee/eDpJE2IxWhwcF1uueh1GtiedNthS7Q0+QsqOPpZn9d+0+Etp5ePhxfgIcnKygaaFg
XesG4gnplUz8tANscsnLCB06vUXMFk6PjXJ48ZKFSVY6sbxB4yDo9RIMCAiEazJ2bOSEQAWV7KXT
ceO20BoA0rL5NAO09F8Bj9F5W4M9WRA8pD3Le/3GhNBoEiSfQBwIoY0UwP3ZkL8d2mATb0WHcmBi
34T5NkFMAyVXC3yegvlI3LRXxZPUaGQ/wz3H5qIvVHKPN3uGWWOL70MLRtDlan43mVkANwkKoNp6
6AlBzUkdAlMqEE8ltiWPLakz+IPFrEs3P8trKM2jGy/WozgcHNOrpAq65Dn0MVL+QqUmC84j1Ec4
1ymBzpjn5YopkYe10HyzkD1cDXe9XR4zZK//E4MD2sSbAh7vPpgnPWWvSS2WCtc+xy4OE/lKGItV
RRHsg8h5ihe8J7c8sqeWyMew3HPlrmozpomCEF/+Nm6ogznNl2wBGVkm9BjZTGh7dAdf/mJPSHho
B1VqVVnDJ5REMMuzUH600gLyESW+u9bE2uBOszGYIi5gT68NpQp+vupgn1dV9w984IMlNinKrjnT
vbszAWCabEh8k07Hp5p0PROCgcAtGa0FHVBDMZHcz6tabkdqK2KRDQnZVOgWRCntsSDp9jGhm25T
utwIL7fW+o6ric4sVutv7h4yY2o47WLX+zgG6ugaUP0dI1DyfSu1mTtF2eMx+9xdnTyk2D4WkNvm
Zamet/BKDl6St5St6nDy1UwTJrP4/z/FFjwsas63TKLwIT547xCVwet0hNNiKpavXxZxKVWppzAb
hQ7Wo6fgG/b2jY+7G1ubaocfJxm5FXXMulnSOiVli02Ofs957BL60YDzJ9LY2TpJf583qjbGs5OH
TmaqabGcsDKV3rCRpWljImRKpAcZnRLTtGZkOFrXwWXBmOWHnR9XfB0CKmAi/Lt7fwKnjpkOjcX5
s7VzT6M27Oq744XDrxqcdKWIgajP3gVQ1H45v+WjWj1n9GZZp5NxqSeA3gKoFtHrgTZy2BZW3nzn
qiguBreqSZfnRaGdtAwz5yosGveEmiW9mrAcCCRH/iYzC0sXnZZGAoaNQgbJQhchYN+97JjDTGIv
T99XAH8D0vc8xkTLgElT0VUqxtvi2zfKRjjIuSolbBFSYeif5JLpLPEw/P0oZnaeXlwRWYzK0Gpa
zilBZZhVLrzory1qaUsWANQ6IPVK4zJCI9axh2zw1GCeiRF00XRrNkna0YJB2m41D5CdTWgAy0bf
fhkQZz63ALJnaLnWJgI7S9prTnCYb70klNwJ0plbQTVmx8MsYMT/3j+iiMf7auyAA8YdEw1UCuu2
QSH6BrMrz16QizWnw5oEktVZyd8W9xENEJn7zXcWoasgZ1DWprrFgLwvWFMWKbg3GJXWD3HeJz52
xvvWe1sgfOvbmN6EtRi2k8Jkip2kp0A5DHCTnpu7QTxFh+hefqkZJhwRQZOqVLVJwIvAHfkSooBq
m4+vUm24tigxuFz2PtGkIDDx4iaqdoBodPGUUUaDCxF3dLFnLy0l2td5OGpfDSM0hgJ226b1cZiP
X2jnXD7mt8927jpAhp92/dVJteYOseKFGtK7P5Bg0FIJNzUGnReE93pSRljeRhVlr1i0UpAYVWAh
a6miTdAF02wLLamHXj4ZykqMBQwpXWH12d1lsUSEoaDQeaWB6eAqrrWqIIAbKRy2WbrBp3ktfdlZ
06jVto+YmWV60NeOcUw1v8vgv/Fkv5nMmt30ri0Pzs6/3YJSVqyOTCEgUbMFO8Iq5J7YCM1G8LL+
zkZx7m0woQN2nrgcXHaN5QnepiyuUavuC05/Kecr6eqj2VsfqBPFmxNpXoBoz8ehGKtqGPPnUMAN
qcKf70RgoJc6c6+90khPDwNF9Qrk1vrA9SZbga8Z+q1dQJFbH8Uzx8U9zQdkf5IPNMVj1EoW4Rf1
IwnUsOchencQTRI/79yJbUfbfcxcJ9j5SS7N3Bem1XvzFEe6g7+mq8WzqEoVsegMIzxfjVqNkh/K
Qb89hcSKGGGBmxutNvpSns3x1XQRCpSbOyQWkdePzZdRlfu7CzTLe8Kf/3KzXpfG1j+Y5eT7L7Jw
ezSHjZm5aUmXg3UYXiS8Nxig3kwZZBcWJJCivcF2V5u9skS4vfastPPSrPNS7fma6GbGJyv1g1td
8Is7byzEe/RFFXUs3+/R71/b+WUa8DYjMUUj0Ao8OmFMWn3u3znqZfDoojYCknmlVztf4I8DIR2m
vtEeijqAo/vP0uSQabSQO8E+HbzkVWCCEtXuQiWFS8HcfRegiCskuviLfyTMSZfZ1pexSJbj5YFm
c5syVbw8L4o0GFA8F/wAWGPxwKbkyLOzUmzbbiV9txmsCrXZnsuaItl0ARS1dOaImZy6R+5uzNP/
98KId3RIQLrcrcL+9Am0ornJU9BjuisMoYts5atKZnNObrq3i7EDB2unPOH7JVj6nY86AE1DEHBV
HoQfJv5rp7uMZKOWBK9lQSRDu9Z+1hRDbXLke73el6iAaE0aLy1G0vRAQi+LYYDHy2MyU+28fsDD
dmCRmWlHDnFNz/baOmGyCutI0qvhnnKk5pl12+uDtJohIExfd0mSf7CDPC+LNdMZlaScsKufK6UW
w22yxHSplNsPfsHsw2UrMSwCSd2KhJFE8dD6FwxcH4C0iimmY1Fgrkfj4R7KmMjB8DogbUcfB5/b
WrTcLCsH0io9bo+00ClyXfq3FpBOG5wuYQ5lgzWoYurka4u0dNRltmydd20Tj5O9lD0jBtLwEvcs
U4yOsPFZmm5+hXWPlNsSyEBo9wbOFLJxDkVsampA2H8KOXm0Inat8nOX7dzBKC46Uf7EkpEq0+fz
Q/nfblt7QmUJBk7V+qURg+TOt4+sdohZL2ircPJl1feOZGZfCNDYGSDq+1Pp6rOJnhKRkM6g3qWn
Pg/wTOr7WdOq1EtCq1pQzm2L165qZH4ipx0EJbRvleKIf7WGhmiJHcsNIqByePJL9ejm/CtCqqaK
SyyXia2TGMOGIhWgeD0VkzKE/MoZgpQybc+D6Q3r5tNBKTEL0LIQdvp2rrZE9WGn9o63Qyrirb0c
URoaiMygJ4kPPubzDXU1m+rb4xUf5TDY49pnggprKIe6zTns+lEMmrCjliZafH94Tm/tWBEM9xtt
YkezYHmHH7Vsj1Ngsd48BXG4qTVCeMvOF5aAV3wesTyPg77Mft9J/j1nBXBircbOSFUchUduhJ0K
lpTxhwOLkBmhwMDdTPv3NiMAv0yEzWtEaov9VUbTt7Sx2UBCrmnTHUs+eGH1ydX3RlkrZSb0j2Pq
tWYwkmD9lz0/Tr/mVHLXedicKeSF05BmV99rkPse4QAtYjwr76W768heTM5yqf6nIcfoskE02zJM
giJicBS+jDyN+q03e4TvqzSbLWrpjyNhp6Yi/OS/zGozjD+eyFL1YtVRJBTdVnXFMYzHIVTNpA72
Frw5T2eSYShkGZsGcFivfd//nNjPJ26FFggXht7DiZD+Xx9QAMaoR2hH3o/7ip5KNxQUwOv2Ig0E
q88VHpme+ClBSfAAfYH6ErBUrn2ymaIsdIx+uTQjoDKZa+d1hqSM8JczOMMgQy2G1uqUXa6AQq76
eDyAdT6Pm8oua0sA122rPU7VJk+gb09+Jb4t6BFG8I1Sa9wjIUTkCnjSteL1snRC+GNrR3+EyxYh
XrWfRZLkhiDIa9tHskM3iN4CEGisbosllXEK8UA++gKtYSddP3qGtmSJM6E8JU5blXF+/6hfGYzA
bQKSdhIauLObop1cdMcqcmBSYjRJG69MVMr3xxbeMYi5u9rhgPHL0CjHXy+eF5kgJpXgSJDyPp5G
QFAtd2dRnj1rtO6qKmCXnaTdyk3mOLTXNwPqn726CfAp25o1puxCbUV9/3PQG8XL5Rug+hw+likj
2jLhax8mhv0HSzmXqWHTDLlY8o9I7u+gszNtLN7EPOAp9CxT0AzQI55lUoZV4kkbmtC4DUq67rVn
6SEjyGYlopZD32tjCwlOzl7IFTopP3mABUR/JwmRuEgtV2lahrg2AgrG9SpaIv2VqYyEGkjuGwtI
6322TB24lkdc8n6xGIM2fja6WfP+BrlA/jSqkXm1Bec0lfTrsQ1H63aeL1I74mEGC4LNZlpSV7hD
szSuJQOifuoataGbVh4vd02lpaG8ZgwgHBJxUBgr+QcZdoz30m4Y2ma/VbAEOj0GzirhohVwdAml
nu1p7EMk9NurXlrPIHmqgB8bCL5sRDd6gqKUHHtRuwKcCmJZHP8ec7IHQp2RzUucpKy1HDOXj+WR
N0rwwSJlndyX1/Z2NuyssobOIK/fcfdwFHuYDxAZkDuR0VA4WweDrUk1d9KL3aI9d1FvLE92TXb+
zf9/XmIAg+8VyTL4aAFvBEKRleXbpXgk+Uh6SAAsNcxVYyA9VJQYwrXcWA1MvfddHVXNRbtpQWyA
S823KsVGbydcoLeZFMGqW0QzdDKQ3ro61ftkXAFt8JmpRVnWV0ECVScZrUB9dMG7UvAnD84Qb6oD
MTpJZSz+tNHkRsd35KNNvWlEOkADA2rnC1OfaSpqrBFpNJ/ENLqaid311PQRagQ3uVuKdw5lU9Bw
tDhASMJOhga8/kXZ8jf7umi6pw4I5dnHuvzx2manf28OeoVwimz9yR1y5kA+g6hpmBHXoOc+DHH5
xUP1lPm45TtOnA84X3EB86Mi4eqGS8bA4zHQWlVxzWR0M5iUOXWahrhnyoZLQBMkzPZXXWgd7HIY
PNPeU3Cr8rfobltwHSnwI70pd4LE+E42pixoWa7CyQbtqp0O9iM+LLoX0n6+cV+EWmRkXL1WqY4n
f+k6pz1nNqRBIqtt/BXrknbgwuA+Yj2rrCU9Q53zTPZygUuLviqOzNGwsPPoedqEK2YcPWiMk5BA
Gz1AxFC8Te1eMmMzYPmhUtMs3ddgSZPzzJoWF/2kdI9yfTFF6oZTNGWX7GadeBfpGdIhiwTnpO5G
mvVaTWTZC81aqr22EPqC/omXQcdLMDV/jLoWCeZwdaahr8Vudno00XuetgkWfEtZWiX4bgJ4pF6b
c3qja9xo/Xmg7bjI6YQ1ajpZ+f0KWBODEoqTLP/TygRofFTTFrA42YZzRybU9QrJWm7y50sKzscM
M1X3bTGQpniyA5F/N9ut7FYw1GakKORGSChv0oA5E2bTgrhl7K4W02o3YU6nqeSdLZQX7eU5R9j9
ckp1Qb/cc0TLx5X5dk7v8xNwCV4ajC1viASyUB/JCRFLURhC4pXqs2kFoPe7x+ntpHJcmYMWqcby
9I8WERbVHYAWI72PZapRGwSzRIVMC/OSMxCkC7MjHqpQ32UDus+v937LlUuzyczPVICaCikHHud5
E4EQkhb7xpye2SXMgofHCs6tnJk9tJ1pCuwp327Iq16KQHaj/MA2h9lV+U+oIOOL/06NOnZ0aw4s
i1PYDXhrmqwlZt3MG7gVylMahNoi2805leOCjXzHGTQalQ3JXEoz/5lhoRsYQHMoHnXXzHzTTV9m
pVPnA9lfSNZ0U3yoitdcKo8buPSkSRvS6oJNnSYfIrixQY/+V9vICnzmKOENoUShrUXLj8Wm499I
nYoQ0Ufj61MNM3wI9qpqGMXJz/1Bp5UQhLrcA1/bZ8jsWAdm+7F2gehTy4F7BATqrYNIPLvHmCmF
Ur9xfN0VrGa/wg2NP+gplouh+nBnmJZtPEcLcKaXIe07p8Jj7a40ORKvUfkZSmfImHipFddBiFUf
mFFijCbFinIVfD14aNlu5CRvR63DJ2MnbJPjgaqszc6UYgG299Y1ztNw/yOnYSkVNIM/NPVhc36T
0woruS4imkD8n84rEtQzJZs796XpgH+k3tb4oWrH/wO3CwyvqWxnBZVjX+gogylS1KPoUbuDjSZO
JysfT1nGplxWh5y/qStRAiguSn+Xwvt0/6M8w6hlZ0xjxuL+Ff22Y7nhMLIyCp0XLbCtDcvLUOzI
XCv+f9CgZgHNjDEq1FTmTj7KmMEpaQLaVJEkmhA1GpTtSsKnI3GWtM3pHIfjlORnztEa2Tbq5xPS
fYJ+eYmZlW4qg2SEvhNZNRGbbQyxO2SdMX39VskARhzbLj9HkxZaMfLOc5I2uj3azHX/Q8KRqHdh
U8zntXSqR3qdfpEoj2NGqWpneVAGCIo1sE9WfhIGmZD10nRkmYl1Tnz221fFYdsysrRc+6vC5uMu
6cAAdmnzXhmrE0+jB3lfH2c1SPoEjh7Tot02UeDi26FEPl/c9SWDWALaMbmbe4nYUnL3E//DGeyL
12b7B0+S+DuBHwKmCAnil215hj6Drlfrhn4yttSL7/8z+4hsvoD6cn+WM4iRi99L4dn7B9LP7Y1c
NgKAHo7fIZ4bSmN309OzoMDzhg/u0QF4ZgX8QlJq8rrkTTrtkW5Tyrf2FGM3BtFB+wRCPfRMm3RV
7Btxgokt1N12qg/LdNppKNGBsOH6Y1r6NGHEO+fg/+fTMHV73Fj9ZyQ73IMGjkoHbl+WAnijtY2B
YnoHTsBbrNWPmNP6cj6rcsELmNVZnA0HUHYSFvIkVzAsa6+HafOjP2f9Zi9G1Eup/5tkkPyVJ9KK
mjFIPtxM5czWb5DA0Lz8MqVMFbTb9xslxFLH0PJY4+puta9rNAAJArOuLB4SSNX4xgWJjLc4jVL5
FSvgBy7mANhg2QScZbiPRPdNC8axyg/18GC6Dmd1DD0MS/MFcRJsl/NSpkXQ4VbnXXkerhh+7UU4
ENqnMsbowqeOQJIuK+oVAavVhxHYaPU9CWVuZwTEXOe+e8yoFxarZVe+Ux1FXl47nFJ1DgCZjaje
MQsCkXgGR+xIRvAYukFJTbFUpTasXw7edeVqt3KZD/lPo+t0ZLwK1y0PGQ9AmJMf3FJi1UeuFO6w
eNtnJlD49baepn1BYcS0Q4LHjdaTZpT53lMAX6S6AzEm1fZkitQqZL5qfuXIPn3gab19j4nARWGG
eOdE0vmc5ff2WfXwaiarNxfwizKbHwf9OvSKkogTdpjhwPJ0NvcPoB/WiIx7eS96jxlBDp9kKkig
mUB2JYSnDr8ccRNqtA9QbgNJE5VG1Wh59H7sTPWpbDmbW0OuW0sfpnEzZ+a+AC643YixJ185eZAB
ElQp4j0b/VmGo2ukz+OhIKTv2ST5R0fzGfrfaD2JDAccVPGXOaCfjyuMc+WNSp/zUIAJc8KG87DO
8zFSpAoC6dJ+aj+xmTJy8QdQSXuQB9U22Dyouh98ul6D52fq3CctscNLwDBGgZRdYi/8maVbQPbE
aLIz4TTAsBpN14afCofB4AE5x4cKqnaF59OV6SFFj68Y4Dt0y8ybd4GRJvNun+8NSy2Xw5gvjgkt
GnzOH5rfUziY+5IpNjtZM+j11xUzpZmbodCOzm+I3vBEklVT+4af0+RczNcmPmobDRfAlGv7IHQj
Kx0PMZgfOsYjdV6fN+/pFvhSuICklhOTMPMWkIWcx8rZ9A/lcr8ZJRyixPYS4Ty57C9dOMc5Hb9m
s1P7nAe/efJ976bQRYdc41kw4iPBJJQBaVp+0QAXKOYcbSP3aFKfPiDPBIKl+QV1pM+kVVfe90YW
dDK72R8uEfHUWIa8I6YJrexktrHXvbZKQPzEn6mg0gUHVEhDMNNS2hsBZlNAS6XN0h8gCaa0VtsD
gSETeis+Mc8Tel+SWbIKxYn7SnUpAbVWgExRznuXg+JTXbVVh2iBV+rhOuu0MHnnDkZQHaG+p71l
PC2wRkHy/i60lC7QAQfLOjbAsWYtJsBxgGZBSpo3RUJX4QuivK1//KkpSgn86xRmNFFZ+z+xgDbL
W3ShzVkSvMGhaapl+BlPYI99zgkGDf7+EzuO7iVCI1v5URimy4JbICamw5cZjgJuVfdDMvOBQZUM
MZoeUaSSTR1gqZeIpJGi0KKqXZIeNliaXT63zXN5wuTlmNhhCYYMsiu91KvhYeGA72fWzBX/hQ==
`protect end_protected
