-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
C60jYPtj3a342ehCeTNORC9eLy32/SPrUAgnb/J9mArPe0Uq1h7riBbtWLiWZbJ33XWfuyVeAsnJ
8Mq1MmPMR2mQxiu8bI9v4n0VM+z8lPz53N7V4tuC45y07JNEBkPjAinh8bDDTE3GqN2vNdvaMRqN
kkeQmLsT5rzjfiqHywS778UwLjrVl+DQfqzyc/ZMlqTYwgtlqiuQLOqwKFdUSvE+VwjxxzIOfjeI
k4qiqZXwDTQNreWKaboFQJ6SlUO3aFw2mZmBn2YhvrORxHb25TZMFY9yqM3G1iWDBuIvPpDmm4Ts
9ZnAVXdeg7FM32cqEkTG0gTRQfdy2V97in6DNQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8336)
`protect data_block
Ct5aYL4ca5m1Ngdbs05o05tlUXtetwVpTtBon0MB82p0wLoANkssJnCrWWwE3kwTHA7S6KxL0GES
Au/WwgCAz+TVATYeZKM1uybslfU5C8IGxy1femW0ikb5WCL2l/Vxw70HUB8qT3BcYbpfiH5RjUEI
8lIs22hH4414HlqZUbiboLKeWcyHsKDs9km/eWSxX4BkCYykAs+Q3R8ERhZP+RX9CN3JrgkOraBZ
A+3B+yy5Wv/3kDf3XjtcoEfy/A3WZC2RLCUTkBcaUA57ey64F0bwn6SXYa8odpu6tJwugpXf99uP
4VGEni3UFJ9nmiv3gZI8g+8yHciADLXpGWc291PwejOzMia5+p0novdhn7Cko0WxsXuaILzagpqd
pyuiYRq4qzb+bhXDVh13a7Z6mS2dMfV6R0pmX+D6KvIyH4aK1t6aCcF6BF/9t53bBmXIfbMMvcr7
AcYusHvjR37fb/CqHCw1suy9Rp8txu2H9GaMLE8aPVK5qaBOuqQW4k0PSs3qpdCqVulKFevvUvTK
4gxaLGCKbNvboCKey8shPKzlHlth/Q/LNl9w2NJoFJfBxCFrGJnnxndjTaZvbw97qd+wZCleOWdN
l2jcceKTfjpDrPefavgvb1+KSTzmoNhYffi10XMQDZKmDA4ZE8bL/yAHLuELsAO8spQN5eSKZPmQ
VIywYG2SnrmrO8kbfjhI6AC/nkV7z2BOyG+EVeuZePozvmSKbria5xysPliErAedXcDMLwC+WwSn
MsDY59S6K0ln9Z/AHIQ2EeZFvKC3Ju1lRgXzofLUaxpXc7h5gkGp1T6CVT9lsIc0MGumhYvBWbF5
lEGKcDFKqDf0IgdlmzL3jh4YPuy5rBmjugHH/goHYBzS7LfTqahysd+Aq6NCsKfFX2xUvZwN41Ek
GK1nzljV9uRutxe3J4mXzXZNRvwQ4zfvYScWR5CD15Tp4/w3LGyx7Mb77ADENqguBdGQ9tnyOXL7
Rqfg/a4tVYijJ22h9KQxRzX+ysVKzVHSvclMKbQT3PcN4xfCJfVwjBjCMK6dv5Q0dCATEq6G3ggE
f+jKh9u2yqoL+Z0BWJ1Wn44DmNlSoLaE9+AedwhHsql2HzXLpiDwZD5/YFM12zmN179Ng++CTGNR
nnx/M0EeH2BiUdDKGSQAsgmklrXuOXhHU+9mXKaUajxiY5Z4hfw+Mhw7XpwIQal3p/g6C9JJbjJa
X0LU7fKgsvYY16ugRy1nh1optr2dTU4XE0Ind7HBBd7NaCdlTPiQR9ewCpDGr8K3HeSYERhkgxO2
e9EdvE/t5gwLsHCN698wANhOg1zVNs4UKEqwanW/Hk3+1v5KUe+7aQxj+O/dqe6VaOZj+sBmZCs7
MKBSrbERf7QXUyFQM8k1NDYLogkp4yycLM2j/GhxaevV9WvOOR6Rfa+NzyndD3kVRynFB3lntcmT
tXAnfiRJMGlelSvNtSfPJs4sWAWceewcb54a75n3I5YZTgLO82RSRHGDrUZuB/j3qN5iMAFBOpsp
werX+dt4G38veiCriseAwLCPv+41rgyKWvuIukN6dEGPSjb4LUfWqe1JeCTmGIDKWZKel1+Gavcu
SaFbiGLkmi9YRXBbYs4ZkwJu0S6bBckJ6Xt4olFbgoQcWHw31VdBlHTkikKCqXI/0w6nGn0w9n2/
AqdCj4vNFWRm6NYKFtcdLCTNxVHMVPF9NbeguUef0bwppHUATGRbr753MDAs6VD6E4XnyQWxih72
bdgyFbc01OeMM7eTGz9C5qgnbe4rirTRQaeKUjKmHAToObUOiCr3FL4HVCPw8J7rq5iRLeVa7K6B
dWbFCrt9al1XhDgD7Smt7d8A5+HU+o/ZILrZprNeG+57wMIDfURNwfi41SbUo+4TIZ8PBqLlMekH
WRnyPqovwQpHHEhB5acDqkCK+T8vEVyaQ190H6BHJaruNL8Q9NTIQye5rZo1xvrpY/mEPuEUzIKA
nnowle0MUUdq5LZgM/bUvEl8VPWdGcs4gyGjBBcu8Cyu0wZaspPNiqf8omwwFoQaKvRyECgEiZCt
qUbGm7QhtXEAHSMHz7haj8TCpZTTf7nJNBiDxXSE9tVHnky/+KPfTJeH6QoC2FnepL7JvAkV9L8O
YQRenI/9j20nB39JSVS/o1i25llUX19+ts/vlzTw2zv19KV18o9pmTt7D1XCdhUiN/tVIAqNhEtz
zC5TPDRKW2iHAOLy5T2A8A47HfDdy1J8ngtxTo06uRHGK6DmY8V9EsIil70WDWQJoJrqmNHiKV7F
btMGK4PZyoC/VHpTMOpujqtrTSfyHHtrKWeRRj/89odxv8+eH4nkxoFbzaIelXToR+a6Ist19Zjp
bggvG80MC2tCLqAi+hWuv+S+pT/Wnu5tQCkjQG/+eWTHS/SWJQhFkej1bnDRzdfZ2qKLRZns11GG
5G90Cakt8v4/s056Aq+flyuPtmdtVGijC8JV0ZozQr+J9XcOnsdnGTjWv7fjBdTX3zrT3pDw9t/Q
i/3PcfkavSex92jM0MWnpJvK5Aq53SnqzIHRSf6FOCRbGBiiyxEwF1k1OgG4VjYyd9N++Qza5R8z
xWOs36MabkBR2G8B+IJYRq4OXy/FFm+U6TCdT3AhZBmLYDkojbDryWsOsmKCF6xfJaXflKrL7uf0
cMSDQ1CXt0x/HOOwtdipq7ucP8CvDV3Lck6I30L+HClXh3uOJj7GVNaH4VFw7/C1dQ+mMKgAWrIE
ZMsXGUcw2v5QeFGbF4+wf4kN3tMu/1H6rX9S/Go3alkXfx8xiOC4m/PXPiRPlXQKxqgRcCNvWqNk
8YNuMjOzHIpX3sunXHqcJTU7w0Ukurd8mqkTQMOIcaDzVl4//kxW95Oeurx6cUNnf9abSqo9/sFT
bq+RJsk290JV0DG5oSf908Y3eMsBtxf/2THXr7mRnPdNtQRzAnVIFkRJscZ5fwZTIbY3dCFLpYjW
dOYUEVXmGjvEk7uxr7EEB7tFOEtfa0U7LL0oBEoyqEMkh6tGYRI24aCQR2CDrMujvJGg7bt8DBnZ
2tx1EQ3qYdVZK4dRvNMBUGEX6PnuZV3Leyu0FhGwYEYSeLl/FA5cEnN15fZ7AbPvfqurcOXoBScn
EvPKuzVrVBPbNXxWAUsg+BqeMQkC4SvxK4v0ZUS6wY4UAv1Vp9u41P9It8pNoQFC3it7OhSXu5sv
V8dQ9vWEtaiAJ1bbGtBNJ3RMLwoc6p28U6XvVSCd8npYZq4cOmvpj1ASmB6TlxCbSQDij6O46flO
aEV+gdiEm4CKeQNv2oE6eNacziPS25paR+w6BcU4XJtfMkKTbNOVXohXCyuGWqj6vMy3ZZrA92gR
PlUj2pqaNX7dKULDnrjxr9lG7vrMn0HgsMrQCmc2wMVKdEudKZgCBRYm2WkJhMUFdhJGHNn6wk79
CFa2cXNGJmqQWny08NbB8m+D5U0Gc9BoUFWU6ZyechUzANGAClOWb0xqbtveGjaHtkVxmHk6hIvm
jrGr+niZoSBPl++3mXZ5CPhb75WERJdw+nzqCPqT5s7bQADiSiEQEJGlf307BMJvE7eyBrk4WqTE
ENzUtajUD7GnlZoElD6s5zpHTOJL70LfOUY6Nc50qkp37mRns5oJpIdNOaDlj3bMdx1iQlA7EANX
nI2boUmVsCLCWmQo0StkG+cmt1xHlxyFV+3GGPpnpQK+cgTSNeDUqY3RBK98MApsXBpSzFjf0cHr
GlpOq9U4zI/AnzGDVP2yEZmMDiP+4+em+dd9JwzCwj7/yYu8xp1q1COM8nlC9p6mAr931cOjTKYh
QW/VGmYDHpSLO2nY7Q8pfM5ZznVom3DT+8MVaNTFc22oIWELw7LCqaBE+PLCipYaS8ekNx/KjzJT
CkY82FZ+XRjpaSmyWiFoIQkum/XIH3UjC/GCHdMgpVnfx1Jja4kfskvQQ2L03uq1k9bEbJWucO/t
24J1PRCAGlo8D/1FecVJc6DFKmZBLP3+/FmK0Xy4z5p60rrgxX+gu9STj6woTCwBngX+gvFOIm7V
CLMscBQZQzhY+KzDNon9SO6iO8wmMB+w8dnJh8InY92Rph7ZocHo4X/1ZoLm44paYvPf2Fv79Tau
QZXL45+pHIP6V4kV3mTzA6pdtO687l+PByXqn7TJu6ynR6eX9MN/gioZR1pMh46WyZHj4G/ImZnl
aU0cwyKZPN+FsBiANX+5nskxGryKuY86N//31J1FfwMvEitQrKIh6h/MzzxNHmSVMJN0Rqy85RqE
WjvwLk+Ow0d5trne9enl9soJluBJDbTb6aCoLFTsl/ouKS85eb1gDxbgXgrqOJWC6Nwf2xE3+tvH
IG3d/9EiVR91pCLpM/JakSbKV5fK4YOzxdbrNcczVo8lst8gDwBcAvwT7SY4YJi65Qd9estNX1Aq
hhxFpZfo6zi2PNj6sktKnMtKGMWOoDWyyu9OheRHKWHdOmUYIgIegAEfXbn2ZLWmYJC+Z1MA3I4v
cSdhi8BgPT2qDe2bi7UGiGcJCbOutqH1l1dZy/Cq/4VQKZds80CkKjOoZcCOGCoqjBM67SYZzWzv
5qbhm3uJaLXmW9QiLEGDVsqtfmvr0vEr9lVrL0X16YTciMiA5TCU2JNf91JbI9eIdJIj49yI2dae
KGHDAeS0ojhnTdHixwquIses7WayK1qeFFRjZuxhEk9rqXlCKwhsSmHM+8M9iwnzrx7CdFnV9BUm
KukDAC46F1WEQvkDUu2fKonS1dLEi1MNAu3lz8izGtryKF1DLYkNdIDx7D4yUQpv6NnruxaaYmYo
QIk8klKnjUG6WAQqk40XbK5By7eowp6AxbKxbbm2poKmvTZw0vRc1ZRPK3pgRxdLe/n6T+K2+Uvy
bBUMbNkeP4743RH7jDr1nxkNnBYJQZP+LTwCDaKngaolabKzG5c/9ODLd2m21AxGO6x0YTE+i9jf
UIRgdxD4ek5xffPEtkvo//2rcXYxQbCzwU4xnPiA9/53hYxKmzLZih7fuk2HmPCw9qnZlGsC7a6T
RGutxmCED5KDGsV9iOrlcUboA4TgRApNaEPRKbV+6Y6vHzSuh54Mm7oDIWxqnWhMSEBlwOvH90ex
LCFo8QYPCxtJ3go0x6Y/zlc283G7lhNA04Eo6xo723J04g+gHvl+EsJWPO8o2ThOMVE7BSaWmFYo
32xvHpQ2qERFoLUK7HPRU4mnIc4bCMpj+63GMrznvu//8f8agoqCSSzNAg8fOgcdyxRfmYHJB5bi
2pSMWBBQ4aHp0ArFjoYlJ986y2gF1iPgBQpxhd3b5v5cIddtEhBK5s4P+pgDSuvlyDsZxwbyPgpH
cSbhDOSqtIrH2u88sYWRzcYPYxm5D6R/98UPR9v/kH9ttadsL1kqeA1X9WKt+wG/mtiXGX81WoN/
TSye2lSAEg4bLXeYmgh0MYDlMSQcx9OXTCww+si0RjPJtxuKtBdElprA+eGIJHZWyZQfaUzm5O/H
epuH5M8mrSZ1Vq0Q85WmBNMzjfiLk+pDGGIh5WFYtwAQshTEiWJ9bVDsZKG/qC+yelkWilN8sGin
rVugVzj67az4INP376xt2UbOUFMsMBjOUVeGXf1vM6CgsMYO2/C6zPtP/b75K6R/PHV2WVFEuZEB
lUFW66oiNnVA/4NAiacKkVCBbrD4ZsShlXdCDLIHWEbsHG6gdrENIsh6796FwrYBrzcHWIDefLCS
ZWuGaF8IJ6hAQORYvKizLwMA2DzX+C7C3apm8bHIGVYYMiYrPhm31ainonySjCswwOuNzfG0pvoF
vE7nWT7ZI30VFk61Tvc+RrRK5TCQ6SEqZRGJSvMqo1GApVurBIjGxQfYNXzmXT1Rx/wKaeZifOH8
wcPvvbio9FA3NJjc76809g7NIK5zzRpkH2vI3qwkL+wuaY3I+QRZ7+NW4L2mYWzbGKUOz3c2Bz0s
uBXnpiBS2DXiLYk5fR2/YY2ncOOTEVssof7pytFxU56ISRTn+u7IK35WstgI+GeY/bqjC7jzuaAw
/iRlww8iD99TmON4cpMVMVCyilvH6GNNK8D/Zjdp82lZV4bVtjcIKir5bFb2w60/OARI9OHKFQFN
ky49b+QeTmTl/iLReij8N9kOV663YsW7qG9VyzoQhsxYzZu/Onj9HcuzHTFdd4lp3Qgb5RYnNvAC
8YgrxPMygft66tyfP73F4XpnKOl//9iI+2LX+i+T8MlsmGBEkSBjkZRDyyIxlTQ7BFir8+PNigiv
DwImK8Pp9tZc83DpYyL8eGziSiIf3Ae6qPMsxa53lAiJ1YfslDjijKhkeauDjuPIc+wfHw9hDy+I
sXhEiRiO636KeTIjl6Na3Lo6KhHuSncZshSEAax0S/X5of42dCA2bD9gdmOkNTdap4G3tvCgIFZ1
S7ryuAS9KGjZbNitnFbwlshEJ4fDSpxa8sBRlJMLsnN997rcS/XEbgRYFdxGRapsipdjtfd49AaW
YJJWAotOfcmEsxc4GQKgRRaTyfF1ckCbau3lOIFvh2TXHb1hikTKnKBbBj/PiFXgCzzQFkgTuExl
ok4ds4dGP0uw1EU4kXwgyPYMA/zh8Rf+692fTXMS1p6O/jDBfQtE/Q2Agv1jiWQH5KyEbKEMTD4b
LgkwQAw1RVV8CFpxjgH0gnmQNEw38uHFDbMWNUI51eehuQ+EOx00WxJQANSoCabMjr/PHOK/nHgr
N6F2lUKzXzcRzl0Dhol1rPUy63841zYctmPbnli5RM2uRByqxi8FTmDRgC9mOX5+vQK5KT182C2Q
sQzAKX8o9j6T9QUsWb7X2EFkBI8ZP9ZOrbX+S9nIMDJV+SZDL4cPsviFXo7qR75/HtOC50Xvu+O4
lRZQj2dae6MT/jEcjZ9Qf5w7wyFca5pxK331Meb1WB0gmFb4aMvI7H+ezhTXQ6aReZs8R6+AoCzZ
SSHRTGnnzdGeEcXkQuxW1YQvSdKumO1GWwaxm/hAtmhUd7mdCLhU4/pSeyv7eaa+eLHMwU5+oAq7
KVT0cOQZynHuQnVQrcDUeJUKjgZ31Tp63uFFbMxw4wpKOZGONuBB67FEHyIoCV4GJcTY1z7i5Yh0
PHyBGzkmTshhCsEi01VbYXNn1rtGdQfAhwwl9TPM8dAu5YL0p+HTf4KA/womOMOaOTqPQrrmwVnd
rxd1qu4wrLn2SURmnqhs6CtzZsCBKeLR4OffoHDtNoViAXIvlu7wZ5czFVaHgC+9/6ws077qowuF
xiLRpdqvEUwmcu/zB/b8YMNcSowxI6Z4jC13NDKhoYZcGWtqHvYEkfb0deCpvKS+pjM3z/7bYBgx
0ydHgdCdpzdIi7o1l8phxg7yVHhm5sEOSoQW6zzueBC44oh3eb+AYV4K5hgHrCyKlF8xvXaQ0BsJ
V4wT/Qp6qYHN8As8MdpZI7rMw2/VdJJM/FZ2zL1jLQ9q7dki3YzfhHAhioMRRynIntOGQr6yPFcc
LA4PB1s/0gh642qnxr8e9Fwq5bcOWb8mnpxKwkX+mGzgWiOQVvbcTT4v+1joYEqreUookKxg+pmN
rf9PC6xJcsDAxXqenirf3HO+NUvSmPo/zJOD5gzg6JH6Zjd+Ku5nhvnD3jGJECOnY0EG4b2Ebj4P
XyPBzmfuoLTdMFmly6xnFLwp4hvbZPW5B3c5xt4VaOiCzn8IAFk+/h8VGcCh8F0kCplYQUuwR/jU
LkD5FpkavcxLiIAW5Dfe+8LVTHEEjxifVQZfFb4MZsYyj5+RK/dw7C0T50mMmVXEYT957r4mh6Dq
acOC6mAlFhGewceEN5zaeNzAcPbY65S5PR5lR1D0xsor7qKbgAjLvoYQ0YWXLjwoSGtS8PGghW2D
e+4krurHmIF5hXQWjXR8IasfZB9SXXgQuT4A/1+ep4ldkjxxN2N/iNTTdZMm01pgN4fmASuoN+ML
XOI+b1uOtTx1yujwjHful1u/Ltto4ehsUuN9hehd3ZwJfOj/wiNlNu6tkJrHkG/sOhtpG/bbRqK3
vSpFxVO5asbUgSdlHXBXLCVNgfR2Reo7eQrWwgGBpfQ6ROOL7/3lxUokC6EElIhGqUF6nNmT82X3
/fJ3dMdCGc+QrXysb+Yv7QS1D0Fb1bWTame37vWhf+Dme4w3ec+BmjGUXsGTfA24RatIGyZNzDSZ
dVM8x2vZxbwncHC/+SfT6TRByDG6nHEe445M7r0J7DvWTTOusMA/BpJiqRmcDnD1ggi/R5M7eVw4
8R9LhGipPbt5WE8KNsE3IIbacC1mU6SSuWyPcKDdrf84nAyQniUt7MO7vtWYP+Kb9tzIjiWILE4K
yARzTD4p6Qc4JBjF/Hv5r80ebtHq588dZvUmJQxftgZJOI4wJfbUBU4/iXQRQsEjVPoFQbCApQdB
Ws+iR0ddx4FtYspETuLiK5q7XnhEG438lwK2rd7CqUcY7I0lW+/HK/Rd092/gohNbKTxzvjqsVvR
nV/a46kEXBCP1m9Iu4Q87ojlzXWDJesbjZRbhepb8E6uy+JM3zVScbviLUd/qnTQvj0dWdC/8qo/
PZcwLGORmqIqtQHC8qKwDlUWygQrtFeY9QFac4NHhiLrr5ZGYbsBylUCRz6y0CKuFkkCE9L/Lza7
IMH1mL/9TJNSFkWjqeIESBxiV3iMAHrO4oZPiAVUSdL+c2f7fy5Jz3OTSTidBlN5M4OEI7OIvn+3
l+BM5H3/ObvgpLqL6uoSmB0eKDmwoXaFEHcuY5Lnd//uMJxZZBODCOEzkJkyHb1O+EmuBChIZe4L
GxacyN3qSfkslS2wajwQMDtUIYhNwxtn5LQKvmky5CyAhFIU3pj7/RkPImQzS/sn3Z0CSv5S9JTI
sZvS0FtqKRzs64hhjIv4eceFB2U1gxPFGgg5sBoZ4GZfKB79VccHRzlCvN/GeKkElQrb4vBWE1Fm
YPBCg9AH/4EWP8+zuUVYiHHoqhyoy/a5as8m7ISpvxgEEptU6lXMLxunfLjFAnIP3XmwIOrNEspH
v7zsNXSYbjEI0ZkUXSAwPRcnWpoqWtRou88OUkWlnywBnSWtBn4tRX+A/HhdR0Fkipb8nO9IeLEH
rBTQQyekWjYWkC6D6I9k92m95m2YneSdsm7PqxypL9EJi1XQpFiE3CvxK5dLQPfeGtd3y5YDoEFO
MzR4uoPq7uEeZKPiTNeUkGIUCF9N2uKh7bCErGo3wSKh1WquSyI+LuvLIjODzbG7GxwbiONM9nej
ePyumwcAnwNC3YYvvNj5IFe4+lIRhMMPsQTfurgIKDscFeB8XVS6hPqermnH/6u9JKomimqYfJjd
N3e8OCy9tzmnosEbtPlf2Z6PE+excqpZQiEqDcc6JwbYb7slPKAp1HhauVWK+KlbAERv4iEvZgd+
xIprc6L0uI+6F/Ei0lNbs3Fa0v57dHuvHUQ98pMfyoqyYgm1i5np/n5NlFtGtiar3wERKepXvnTk
aSNXAbRB7j3CtYaaKuQxXuAqul8v7UcAPhlslbVa0pL1WuSB2coQz82w8leJvWdTPvg2ah86XsGV
0feC/tx0+A7om5Oan7xQXGN1kpnQZrazxVRBap5LspbR8HJCrTjheu1h8K2hzTQb9Y0fg+qIbWDW
piSAo2GttXDcuDYjkfDwDJ8NzCfWbqy8zNW/ps0gm1eenJ7yjaHKYNy/XGkCaomj83NrDAP2YtZl
8SZH+5lQQpeMOkvW/Brt391ZsgTyzdp8VYO8CWbplamDR/+81Mw61sK1YtTpoj7mWAcrhKZONY5E
4ErmCbts1Ng+boevYiZMDRq1io3D3lM7sCkjKFMtuwl/6tJYENXTZdRhy8s/l5ArD1my0gbs2uC4
XNh8MxBxA0rwHopPv9Ydw+V2qbzT7Yn8v5b7Zr7LbblkAizs+brOasnkGuRjG/D14XTUmKFXcH1H
v6/BSZ6PCJKbT5QvH0zj46kcNlvzg0nSCI8CakEbhI4Jj/MBZtLwGmVodaDowAbE7NAqJcpjfVZz
96ShAd99pwobaw9x9eMNqCPhtjlg3s4h1TiyeiBPWYKfwUhqsb66gTzoDvo/RgaSXX2fMb8AIQjl
tOlehzSJpM5SwtrlCC67U2RutYVeDEMVUig0rDUFRBvvSbSwI9C/9t1JgIDozI8OBJOmufQRyfZy
aClg18+U9ZUZljhpFNPIQXYYu9gZhYJ4Zm2iJA17gso77rxPUaW/p4Fs/QQejVYDeMJ7lczWr5iZ
WfDi5dRv1fygjcfUKOx+9+b5LnAxnVj9QmVoySaT/tBXdfG17tH6hlwQlbuNfC8pLyP3GKZAZBSh
UWhyvqAfQeAiGQkbaakhjGBYwo6/5G+bbO9Je4E0oZLVIbhCZmO2QEaozMIaZcjpShPhphOtztNt
vafmQJ1IPLknFXhrT05+fyEWwTXkr6zi8ScZzaCiLqmSwGXHC0+Cn8PE9pRkO8wSKupOOAxCniB+
yMedWCnBM48p+3LqjpmOIxhsCs27hYIrJvDlrNQrk8G8XXg+f9Csg97+G6mYJdXSTDLdpdQrF7LJ
H4vbFdfyRGzKTS+xerLJkHG4XpBzYmvMXXDFfPxkagksT3+si1uT4dhYv6waHe5NnqKWDLzswa7+
A76fC91vedKvSqWWW3WjpwbE69OId/xA/zFbe2lbD4HBdN5ekM+WAzF0oDO4E3+wMcT2ehdXkUnC
WDQHwkZJ3+z/hJymulrKyvqM9NxikbwdDkH37akttifan8U7SLhSaYBSxpuvFegw7ztRDCPd3P3m
VxbbQuldA5vWrRwChPiMTcKPM7Td+v0trmtHJ7L3Lo/TQ8ggcueRbnXq7rmjV8fmXf7xgkStUE28
/0N6/OMrWMNgKkcVEyPNEblmBNBopAUo/faf435MuynMofJh/z7vvhoidF3kfNaY7vSKDQbS6gzP
NhIpRa7sDX9IdhDbQCACYovYv6s73e+1hzpq+uwgiWkjSgzd3M981XlYAd2+UETBAYEiWjUXWljz
wRjh6iaLuOMvfcp9ruwvy2elrMXge2yGz7ZXoyI+9fMv0tbOrPsV4zJhO0U7Nr8uZoXy4LIXNQto
RKsGFSvOcWrfPt3xyU0WlOxfo4ZJ0KBlNaeBsibH/+zyWusF+pxdHuQaVx23cZ/Wyi+9YwbwdeEc
iaVxYtqFErKTxLwDg2A=
`protect end_protected
