// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Sun Sep 22 20:49:28 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XyiQ/QarHBdcfDOPaHUKdrI1pXqbVtZ5ZZjVhGdjrzyBvIbrRizzoPNe6IutoqBy
7ZsbsHxILBX3PvbiVWoi68nuNBBcIOjaguv7x5AhU7CpFzhdcaYcLMLUFsto6FJD
i1Sia7w3Ne6hMdFkMcm6ECxZ5vmrgqCNxEiY73OiDis=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20624)
6QHbDGg56/VPxQghP+UHAaJb8c5NnNq4bbYkzTotaz7vful1xMCpysrxgWiChKIG
T1nvD8J7XQtlWdUsDjHQjdmOYWYn6uCjW5OUhUt4j0UqECX7ag7R/uX4YmYZgpku
Swu/PKhqxnqvdpLnn81liX0lc67E1R49RwN6BwiqidHRoSaYaYC6a39/12sCYF9W
jGztMXkuQle3N6TqYQBKERYyNn0rrOo5RBNyVYjGPkCeJ53LZTyw+S/PYjpEiSGt
ram8n9nMHv/efb+odBBNQat/TBeOgDnqOnGkLH7D6qnm7J+WdJld8h6sw/BdsyaN
u4QlUpCTJ92m56m5qXCQwywcLmZoBwrQ5qn1GF9bjCnui9vjbJJdL4ZNxQPv2aKG
AELpOE7ZScsIO+AElaKIq1TGBVBB/QI4Z1EfY978V/618W0ZQHxC0IGZC5y0zyRz
NUUS5NGut8HMpMmafWiGY0H5wIln4+7cB1JjL/f4WlGRan0fl6exenfI6eBisAbr
8d4hZp+5ywmWADT52vmfx4GpY8Nil6vYpBO/aHytMG2F/kqHeZEdpjpJd6KfWMTp
SrIF97NA1zDeII66jLcmroOntP5Gu4A9kZBUpcMoDy47+We7hYYO/vd8MedXkEiu
RcAGXjpP13DMc0pQ4K1ZibwDsLkkNKwJwDjDdt1vBKyW/nHv46w3WglaGPZ2D44V
/xkb35dGXogCQfQryhFODfmqPw1fvz3AFf1I6wQ/jOv9OAKnW/XnFGEKv61fR8VU
Jt91sB86x5dATORiMqiZe9Pgn3DIauqnUIep+KBXi5FSi3n8BCLtE0XatYaH/vYh
7yXNP8k33GOK4edVNc5l5rKj4i7CF3W7hanUUverAtRFrmWC/N0bZPdtVaXEo0cF
JulOPGM0VCvBN1zh1WlYUJU2Vf9SRMY4Qg4zsdMobQpDmYkVfn3Q0BZmS1P2aI8D
pVtboQ4BP2PDnkvcbFpfqk4PHdftdjEfgXq5Rj52xLsQabevj4nQH34jCrcNMVfV
shTsHA5LnrWJoasHH5CBTneqy/kovGPzB6JNn7g18PwtZtnJOfv+IYp5asQWZ23U
it2XZHw5llEFhp8aWYgY4Rriy6XY2VhKQ8kib/tcQegCyXhe0qVOYRX+mQkYZBo0
vjZxoSlzJZXRYu0qiHpKfqT9zIS+l2Rpyvp8aHljCWBDJlol0bI0fTnjxXcDsVj1
Grz83ZgQvp9HleoP/KdJRf7zognh6yGRhxyJfQguf2PB7Iv9yVqJcHYagWfVTGkH
BIJQ1Jxm3dOZ3HnsdYSvgJXGbMdNiB4mFFagZMl4IBqUw/EM60O43WH6CRcEIbNl
g4ynNYQZmsv6yrlNKVia1/VH5oAZNbVwGCqEswhTeGRtkZcMZ1iXQKA2MTYXdx6V
hi0BKA35aPinevhlKgX4bTwubKp2gthJtbi/3U7+DL7hwcD3TxcmWfEgrBtPwnfS
i2DlCLTyV58tIvPt3GJme6KWkoixL01HIHm69LCu0lUPXlC8E7/84AePlkOr8rd4
eedVcaDU/XXgyZgHs63cuw8jVw5RJFpORTAPCEzbIyQQdrZtdT9KCyazRr9ZoAIG
r4a0JDF8+MYL+BfcSY9SK3KXDr8AfKpsJ5DF/sjFrnfj2iFcawop53GgyjhNeYul
j4eK7rnA0/ki/ZKCqK7/PF5DrdUH7frT6+S/OTGwor8Xm9gFhspR4t8in5N0gc2y
zcuGINMeCQVbauvERXBMihs0Ip5MiFy+4Quzv+mwNqPN2GGdq6MtJhGKQpvIDUU5
6OKTTjVjdKDKU0Q80+dxyKsxR+y2y515cnvUKa5sC4uqa8EQM/19lWF0pAvJeyYC
bS1TWhyYbQtr+fI+atPe74zcMRLFojPXjBMLmZMhfBxFu/RWcmgm9ka89yRJLhSz
YwOgVW/vnJnE0cdoFvuW5n6T3lcCQPG3xNUCBRHT4bgMhIORUMiTBs7YeMQBMVou
Lr5kDza2dqXCibFTQbONyPP7kMa/wEUgMMiu7nRBzn1y9tUN0lYOY0XEfUqCeEO+
5Mfee4aSSNZOYA7FQCUryjHH77A10m/LSzwcqgdkb2eeEdxlBEOhIb6l+XBxxbLv
WDTm6gXm5BYhk/oDI6N7y1ObQfQnYazrQ+u7x0TLc5xXNqx9mAd5JMnOJS+/ZbRX
QtwV9Zqk3BYNGbuKhjlPXsNFwiORFTao4LN4EmJqmAYL1QdIjtG6rOLqjX9/1tOs
WnKrKUxEHLi52jiQZX39Nz2st7tPEzRrQa3Z5dFora2h1rkBX9qsYeSl4bUkyzD5
78NAm2UHm8ztIORnZxhPDAUBiMXehYCAwW442eXybk1YG/XW+IVY0ZLXsVpce7mk
vxLs2IuEYfMQY+PiRNdMtxn3KZxbODaoanR3fTM6le5m0cXE0Iw3LVBI4XIG0vMJ
lW+hIaCe536UHAvB50BFtVkyuJk7H1A8OzCjXD27Mxd3D/btuj2qcOmWEL5QRjDC
X/Z9hkQVLJcspoVDCnkCaytRdcBNrI0JcLWQe2l/5p3NdWE5IWpqiNZGMhD8p/Qe
1WAXWoVQcgBNabennttYOJIjYbObFuWrAe5CTs3q6xFdEH1ob8z8kvELt6YDs8Np
3vTXl8gXln7Vf3O150huDerUpnOmWul2kjasiTWxUmWHhxT24A9Oxhprwh6LHL5A
lOPUMq7+iOorD+nLRr3QCrris1fYMC80FMk10QwW2X/xMnGtHKHHek9pU9xgP6H8
h0xe9GMY91NWv7lqXDrNri5V/Ogsp4DfRXQNg2h/TEYZYLNB8KHWDBmnr75xbRk8
JZMc4okRUiEGNPMU25M6D/xzFaXTJWBf7NrKZrSYpvrNZEvGB2LAr+kqoWnCUxhv
Hc/1oRV1wZLBEzXKrwFzuaKnz6WiqwkfpeTQ8lGjNrBv039ISHDQbkooWPQWYUhH
UM8qSjG8XCe+u9HJHf9ex0GP7m6c1DTMLwBlLvYWEUu0XTynAWQuWMqXYpzvLtS3
BUtKO7P/DYviC9ubeih6PNgXg8PaPk9BgN5oAm0OrjH2O4nn3DLNuKKF57U5p3iO
Uh9gAL6GYSdUGzsXEOdKyZpj4KN1RX0Kp8W+24xUYfJdktsgHelnSbj8JP3z5nGt
GigdYt8oJnaybMaRGW9lNR5WEtThUc7L2lRvVq2iOu3uajU+twVpfBCmW4cwz/cN
RSwuCAMrruIN8nx/Fkc3zWtrCywdsaBAOwqQGnFJoqCqDtCCjWSyvN6Xeh7RDJfM
OOYFxoPGuvuXWaWzW5IKnQukW152zDb9f4SDpM768zutJjTQQpNrGIN3BqTO9RAX
JKVmD42vrpaNSOVObmRQfO6xtgOpb+HKbx8/msp1OPRKP9dhJH1kiaCY3Cz735KZ
2ViogopJEylEbgjaPWMbCQ86zVeLlboHUPgpUtChCX9gMAtkYvRR0o9PFS0G72Tu
U1Fiod2KpmrhZ8Up3d3xk/vkinaK4hQDuQZEHjqj7izEt/nIemgfpkwgpKweKOXv
KymhyHqm/9m5vou/kzt+QcCBWrFPpj+o5kc+x4i2VLF9sm/AczdY42z1J5dWKd0Y
UejoyIvsQq+YwVqyKD3mfshoyPJehl+8c2jE/R9ks+vGgG2sSWeV7100rDJ9UIwE
R0iiP/jOczVSU2N2cFEl6FMdtHEt3XeOTNQu/YWHUSDzTCyHYle5rydG+pUDMGzP
RZyuKpckgEQRRSUtyq1N61odJ9xomYMSRZzjDIThOYICZIPWbzbf2sCTNoDtgBv4
kYscdTUMN+H/vpuTf4m3WP0/Hm1t4/R15cRPbBEohdjk/uW9sB0yiXB+jMm1DRox
vFHbn2pKTRg5iGPUVdQ1LpH20OHa0aP0lGHBPc/ard3y2BJBg69VIJVvs0E+cBzd
pyklFZgTqGPFQxeIeKCb8Kj0J5yXcSlyrlcl7TTXGqWPnzyiT7swXpsRPemlorZd
9M28nyqxDFihTFISvw6P5sO73e0j1gZYR7x+bdVgwPLlby4K4WZPW2Mqav9/+B6P
nNhjWYHCJOpu85Nn0hxTzYWtXB17xmUipuUjQ1+u6vYV5IwNC73SPr+HI9vZhGeW
5vQibu/JKQYGsdU6kJ7/6udsoWadyez/KFUTHjojHJGZlUkgecqgnigiHYqRveUw
BNKucH+9apRxJon8xhjKnATau8R3Tacje52VkChcffWtEO1IjQzVTESne1SDqWPW
U0qJhSdQDT7saXEBJJApuIhSW/a36qt0xrxiPIXxXOBwoxf7Wtrnqg40BUC6bIIB
/ox3Zboz/Ha88wQJoxYSZIzlS0DsxCjGqomJ/K/pgJ80S94p6Ij0TFhrao+LEOwi
NSHNeggwbVRvMoUNLkwCGFdT5sFC5DTfDGsZ3d1chTmLkz8Q5YeHAeArTZFAqvte
/6hTYr3M0pRizgLzE50c35uIIPwiPNCvV1S22nfUeb9eMUmMx6TkPeWwqMwMgYJq
lIZ9WnosK+8A8cL4L3SF7nAEl3+zFpqua16NbMt7gOvzGuZel3Xg/lX/xj2Ab98p
HLtprIObL6hpj9s/O/hHA7Ilv2EfDGid5FCcx7he4cHBIrr7lo1huD2zTtuZrDtV
wKWZbheyKTNt0s6pqR9+g9YkXZLnKuEhPVuvxZ8kqmcyvum7Nvt7NyUpyneZCS5J
EKI33iL3JP1CAJoPbQ6dw4vVt4qMZ6CKaYJA9ODZH4vi0ksxm+UMwyZpLGJf3eVZ
l3ciHxfnBpPvOx2G9p947hpsP+BakwGyew+Q7akgendMnl/K6ETLzfaLkFppOcCF
FqB4JgDa8XwaCxuTpBwFywsTNl0SkPub/5UnAfQNFoiBNvM8o75YB7L7/iACjHjf
Gk1MSWKKySoOKfwlv2JP02C4SvPhDOznTbnSwoG03wJvzoX+hv+A9MMRw7mrBrft
+Y03b1NVvoBgbGQncQkAKJ7EAPJZ6tnIqNg7vD2yJbzWpwIaErI8wkoLdaSYXnq6
NcmZhse1Fx9qePjj5dNJvTYU9oHCKjna2rpqquVBysOyjs8T4drN6X53ktyc96Jn
Rl9LTyh3bgJ9Q651i6I4bNGnUDs07/0tQohDXitYnE6TpPKc19bBdQiR0Hv/OScW
GIGU27celLtgQDyCATE9nQID/jPnt/qxsxoj+IPgDVKJh0Ovv+EDN/ACPqSLghVo
tfwWfnRxXQA60HXi93TQlntm89u0hWIGnMAdAYS7RPdQr4pnSAYTzhXor8tGsuQ7
ZGmQwWFTgCnmyVeXCt5GvvEBXNUKGwnThHgGS/3hkUyj16zF0Hiua27ZqGW2Iw8H
Qt7zggA/XwwUCzdNJ8EOBNiLO2vRhktzDq1xUOoIeL/l1aMgH9afSwMYDusgANn6
0rSqpx9XnS1Un652I5czUbyF5+ZfbOdB2eFvR017YYIeR3Q3bXPy0z+MLMaaetRl
mDLpYqeY2gCzL7ykR9a+odCgrJfdFie+Koow3VW06YBs04c2ttetjx7V6hmtCmwn
g3lW0XWDCJ8doksFOelTELboi+ZAScAGCWEz9xcI+YTP/xqVfVliZ6lbgGP7jwtP
lR/1I+sRe4acWgC5qIO11DSAvGmCE5RMfjoZabpnXU0GAxbeNcZEyM5mN9QPE3cH
WlC2thxhQZwPUcXmDsh3Ue5yxcaryukOZxrTIavaf5XPVLCaXeD0pU5X/NAWWXc+
EtKUQNiYFbIz5E/+w5GXXJJ18f+aDvETU4gZd8r0h+M5w3TY0p6PA5J9pP6ShjoN
XOpDBpqp0UHV4K21s7YCcQ1tMgQQ3+9kRJKYe9XrRkMkr7KmjZ+kLD/pB2/qsZtZ
agZA6cHOUovc7ixS+wL5tEL+wU1eG25gFuEhrZDrJE6rIaiaYI/B04fF6UuqZ9O1
xsXfKWXt+TdmOgRxzYQgAPrSKn0V8J8YAUG/LRts10BUkhtkQT6Y2E1EPRsgfU5C
DnxYmNvcETM56G+lSE3r6HOjxWO6KmJG3tTAV4bc+bMSPKErLejfaLVxNtYVsT/l
0knbDQYpeB3OddhYwabAQ92rc8UaEKO9imsAtpiW3bHbWWXufgYgoofuA4vb4R3P
iHiHr+HHBJ3613I3j5vTNaEnIgO0gzhn4J9gheneQkqnGckmuY4CqWj2IfrPX7tP
YFiCikLq3pfLil6O6Ymp1JydrkPdDGqvtWb5xjj1xALjpcPs/kLmZPARpVgTz11F
FABM+i+oSFZGC6mdaDgdFtgbUB60bEQzXukfiWIlKgUe0I0reSn6zpL9pzo6I6Eu
E62YF3xU8/Xsg0n6XmJHwBl5uqrONIR+FQtlKSCfCw7liJ9zFwbUEqSEaUWodlOq
XvSJcDDSlkGqhY7Bgdy3jbisneX8Hv9SsCdDGWvd7GG6+mUT0NGYFXnl6jphmEAY
L6hD0Oq2F/RZWuum5VdLVUpHw3jPuppAV95mmCcbApKw70ITU1a2oT1tjv6AVM89
N0D6F61nbZOmxeQX4yvWsLwewdQSs0nk7r72E2a/mHBYGianJm7wrMgmDYidU+Yy
7a4Wwwf4k3GfSOcL8+70uWvdQw0A52j2jf5Cc4LFHQF2WHb9fTIMziez2V0Hzl7Q
7MeaIZO/lSGNpOjYx1ZL+DfPvsE64byxZTMFgC99Ep6VoXDj8ulzV1lV0u8HyWMv
Q+trmT1D/Qvoij3Y+9zw8x8y1xhHTXIYYHlHwtlbjp8I4CPoIEDWzYVoGULcK+8c
Zaad91Q4wyI9EmIU4F1/CEfl7d7GtGkU++VVuFvuAESZfSC7Ukhpa8PTPLFkUCFu
Pycld163sSuQ43pIBhI21iuMvMj8geqReqD1plA7RkccuZ2y16FDynIo/PWTB+rN
aGnKzhT1DUOq/7trBWyVtoYw0EiK39vSDkFT1npG4cOC1JjBXj9eP73uUvUCNYUv
caoWsYRgtpmAiE41TI+AuN0rXO5OO97ycngmA/fxypmPSVPVqrjw4+amWXmIWyG7
GlJ3nuOzmLX5hdGbpr/VVjsU7ci26VkDVobojf25WAcpxwTk3yzQb/FjwifT2XiZ
8XJkodCDArP7Jp8M731h4XpQsrOaEU3iIO6nD0mSq+Qu8i7s/0PFXQ0Kc5jIZCd/
KN8HQ6K+yS2lHNgCm+aH1lFf7g9loRrxtUBZmXpdWcFE5Odx1/NRuxif1/epUn+3
OHbvj389Z0FKZw3NnjWal9QAzB7XL+Dedcth4fc05A9mkczsQrO6wCOhBkq7VkqV
WC+acDLWaBGFLSrQFavQ6uDAtX62OHEV31CfnYEoDtIWvR7ilfF+8xa4r6Tuw4kF
DaCEV6k1cWjt7aMm4q5P3z40jyjCLoIPlLV+Sm6ab7xCqixypB+HWKuFeRV18seO
SH8I/hKFcGYWuIcKmudXGfNtod1pE1VnkB+SJ+LXyT9cHLRESHuUYbcDhxzbvjyo
jLu/sSmAA8XBP0k07w6P5GlOj8OxTWHJE9BR0ILV1cXRsuewfTuMR15AstePiu7P
EsXuyRZ68+Z8W5ZPmKmGLVB3HV7xMW1o5vv4hnodcF6nIyMkNkWyzWQhvMm5OV5g
SFvkZnW2zDxYNp0yuzrJk6pYTvz7w9xKg3Hqxg2M69PAViT9esK1kZ+bFYhZHkj5
uYHQhyTvUjSppJo0dR+xFQmwUed9Vx2GDYH3/Mm4V6zmTdeR41O4YaKSpsvoqzjT
h66BBLvovFdP1KZ6au4Z8dN5ET8PkTwznCMGmjW/6O8vpM2mRoYVtjnoodFvGJrt
eP3G8S7dl7jwKdc7I1GWnZxK39Z23jRHUbtLO2UFqugq9pUtrT8j7hg937fe5sxM
6Uhi81pjJdIWkYjnf9iWxLMp2+BMhSbd6JRqGSXz2eH9KLQKsC3F2dssPC9+Lu84
IRewB5mSDvTG4pFwyvKI69kYtQA8MXsBb6K2dazTnSJHl0Paee3NDRwXjRkbwK/7
HfVxnBAcODQ+eByXXfTTU7Dd/TtaRw3kOoe+YV1TnfOTHoOuDJH+Bvmbz20dLdCs
AvP27pj27RomEwhQ5QH92myz4eQtk5xc/9cp3Itr4MqmaIppTKF1Jg/q96GzAh/1
nqykp1KEP/Fsa5ZdawIwYzGrMztKSuqPTvOtY+vfQMyvC3h6QiOcWtExuXugyrTF
5HPQd76/+YXvbu8HzltMp0Jy3KflsJ5cDMr03mDUIKntNfKhqBCheifQjLrORo+v
mPdCjt7hv08FIi/oeiKJRjVFl2RHBFwdYo0XF6TCH9JAfbEcCvHCh7C/bYtoBe3H
QsEz4EjUB8Ek9ygcmN5hEjrWvwbISWF+THL4gDHYElWgvt/J/TJry+HVrOsealnk
mZKPPLokLQLT7hQxCVSA2PULbRMbX/A3nGhCiZkWXP3sXW0lQBshJ2jo6l15JqnF
FntBsVFMeF5G7VqJCud+DAJv62fSjK+fZ0PYEMALbHmQMqrnp/2KXk5+ahZWDC/w
6lzB99uzWRSq+QXMNH4grHR6E8r8zvudfZnzGz/OijmlSm+FgQaHXd4lTCXSN89F
3GjTeG/B2DTALEs3Uv1+CMOZvUXNaOsNeVOOg2spM9caIe9+DzSGnz4i+cW/74/S
StuIQN/o7mw358DoqoH1J1dNI+ygIVvi7LM7Cx2Y2+mo95vjlkerCryZo7SapQW/
j7BnHk17DIb6sxXsJZMDbvIjnVYMs5RGOE16TNFHt9vitGmljPKTSiCYbb4f27Vl
7qs997bBCN3Wtlcw+MsZD+XpfUlZIVcQiNoRjUIFEz/ownT2eRE/jeNxeVvdkogE
eNEz01c/hnKhhEJZJ28vIdKdnPXaMgNeWhsA3QjM1F8xLmubdGSt3J2NrpMJepLU
38fVtZEfWAossidgoDdD8Szs556PPFmQnwW0ooEDlvERo+T4NAuqcFocU/spHeOI
N0Dz8T4LP2JdJ4MG9BVKxDTxgXmMLU7Oupv5CvOR+80SAE03E3LIqj5jH/fP8n+B
3NUfiKfBGZNLnz91hI8r+Zt92XXIxkJ+7miOj8GGzQFhSfXpmRecnTgFcPDwu5TT
GCoqSw2qjZ+6XjNyenQRJgf6TwhXnN7ljQd4rXXHwjYlQSQivaVTt7WEhaUNuzjx
6me9zY32DPcSnccjjGcRlWjICyHoqMNevlXwc/DtGnh1tUYSawFT1USO0nvhXUv/
DCuUhCeACeSSXuHEPcM9IqZM66mmRspODVVuYODrP0GSDfTgrbOZPEdhfbDrQL7d
oYUqXWx67NnKgBsUlH5lWTFkRZxEEcdW5ffnlFpPPKK/0knLw+UEjHeI/EoqUshu
qO3EEjepdxD4LBx4+sMDR9BuWvvm5Ze8jFZnkjGbDGhZow0rxgqpu65xk+NbGX5X
TV3F2zYx3VKvbAWdGmskk3i/FuMNiO/iT86SZvZpS5P/ReuNl0ka3zSERb/RZqD3
6qE7EJYqbXZTYf0apNbLwWfbtVAG95Vxo4/02mj11n4QuJ/VUnAo/4sHvZnOypYT
88X5A0HrFz6FuGxq3p7ScocSFyWxz4E+9OXtEoG9SsLo1e8qNJOe78AhL2lfhUJV
R/GNdvc5mDatN0J18NJ/QePUZk1s/6gn53iMdXIsEZXGARrW4sMNuX3qZA000Q8Z
3oDs5ZtGmDoCV+YqWBfO2ozrZ1QM/JM2wzbFD95jasxpFx4Vccl5KGgQHwzEMT7N
lTnPt8XPiD+O1cgK+/JtsDUwyZcHn7oolAm9R5Qbvys+qZZcz1wKKVFTQF7leixU
MLLBwcENPRp708VKNSHWroglZEC7Wj1jeDOE+LPw1AFIBjR9x58aLSSPmCVm7Ig/
BrS7iklX4J8Rs8Ewu4KevmwbgJC9qXmnutP0/9hqeqnpa+V0TAB3/ObpPxnCRlc8
Znq4uT5gPEhWh8N/woFHjPnlXlAxQfrIvWbXfToM6sSu5a16c9B6QXYVXNYf0iCS
o8SKsY0nq7KX9V9zZpFELT/M6hH930PmtNy/iOUbaDEoVY7gNNNGCGjtJRHyvRMN
tEFpP3LbI3G1JRHNY9OkSVI1JMA4lWD1vVPexfkczUHrhrTZeammqY09kq6gic6C
H+a/RGWVBFa3RrmWE396hqQh0M9KXL6RZDrmGxNGFCGF/RHrBxu0vvrzLskcuuYH
EpF7LmK7xkgBEqSdGBxrSv0C5NJMPTMPZJZzelejbpOhvc3ypJOrmBg6GV5QyceK
8lg12NBaZIUmKi+Ec681Dna7JX50iaMH7RbaeUnXB8FuKk+/50VZEoHWHX3M1SSi
8rpwRA3OvcH3KZ0/mDAN+NWATUGomJpl/KQIKwEuNWLPdNlEh6BdHtvuiEuw9TEX
jXH1Gjh5e6jLSoXRpQkW6GLOthkwCxx4+gn/z7gs1n6EErVL4PGGS3RsRRmIDg1D
Sp0o8CDSReOp0t71ebUv47T5HW1bZCuJ1EoEotHS0vycWIHTcGmjFWn/OaT+dl9Z
GEOLDwHiwXEIUp5hwMu+ex+8mYfvm3uNj/BNlRkffw8iCtqbsyK5TD5jJszFoVms
lhl0Go/owwnWVJ3REaSDDuT3W0IlUnMgKZOPnMar8Xy4r7PM9KYEHT2hMae053z0
1Yj+exd8D+3JP7u7z4MHhgIbUnJ+WEOAZTDMd6TbJ52N5mvcOEJoJVaXOmk3wNHB
TpvlSWyoCkVJ4H8dGrKkoBZ13EJ5Q2dzqVmimFN9juwJXzWkqOztiUbs6pBJf3QU
eUhcvI9wuW6TdnTv18J2Xg2C7E3kMOrJ1MhpnyckWSGdYTz9GzAOnsEsujB/E0Mj
4mDBQQ+jBqCkWL4K5E/ASRPl4B6nXTy2NRvb9uOMRz+SqfCUze1ljjrZ7hc1MSMR
csDdWbF3fHOZ2L3EO1tKkohDQMIRgVfZrgbafOR9ormlhCXHk6n21GUn87Z1S+3F
owCq7vpAVaF4G3btbF+G4NjZyxiKCWazCx4rHKEpH77zy2TGQXdSH2uEgQEWLzj4
UvbjuHhJGLPbM2lDefdCi0frsFd++e8JM90V//QCCTRRMQQCsu+/XcDVMxPBHFsY
yvD5rpGecID6SAEEMezKpTc0/xoRRKDjT8ceNxOoHZfR9OMnwXe9CoHWSV+CBtaa
QvTnM760Qhp/dHrOj4vaTUqQG15erCBPmiAqnDexOxV6UeqxGjZLkNW3Bgovm5T1
WOX8UA/latLrdHUPCL3O6qvmqfyqtcG9hni8XjJTSRsXfqVV/D+utaU/u+09BFiS
Wx+VuCejgHhZ6t45oN8cUHE+tDqqhAY+Y0yRAwyj8T831X1GVP5nZBh2sQVaJrqj
u1v1xdJd4NNF2i2fgDWwdu8rTib1/NBG5guWyfQC7U63uvGbVJSzUNx/fRBnRlzM
yuBFLMyM3Y/ClB5CpbfOircyiL0U6hDjFmLs38BCm7xSqfl0TO3X+hfktILQhBz6
Kfny07vEndVztlAsW+gdDVfjMkPlLM/MBuYNEw4hLa1kmOj3MtEV6gIeJPfsSSAA
+52RLhwmgwpaoUOKjDd2HS1BnyTOk1MuacjUUP7T/Ewrmd8M7dO3lQ0VzQQ9RkjT
V1dMyv0udQXpwfSfEPT9Blud65PFOxtxYy6eHZYAaKqjL3EGIZfGtZa0vQvjkALw
dNfw4wLyXyxPwYXiVqXBkzrhtdJvS0vLkqnwgUkLrCq7jZcxCFBP5HEybX790RNd
1olKuJJpNJ8ExRl5CfbDVmTxPx0IgE7ny0bTaHX1MTF+WcLWeOvxLa/nKCK3W5FF
5I/cqu8Vb/hme2fenSX28OrryoR5c8NFXlK2747CKGfnPXh77RDj8hoJ65VFX/QP
97tozB88U58ZAWGKbOcSGEevjgN35sDrv0VL7ub7v2ca6YsSSdBBJKePndDvK34Q
zab2+oQBcee7A+ng5SgGQz7cQ/7mxire/QBG7VUadE8N4IpYy+ss1a+/QUKp+fqA
j54JdKdgSHZ9eLMS8uVC/9x+vUYE3d3Xn9tZo70Hq7nVeAvv78m1B7JdKZbtkVdc
S34JqV/U7OWU11qzpDVyV/TkXV9gisdZDAyqhxpT02XvC7BAcsjL84iUe+ZJXFTU
hMQCSy4CigMVopgBeNWT5Oh4Q7GwaHtH5bMVFE/7uNhS2mZhLQx3o+/DzlfMn0ED
/Pslo1ata4WhHBYZ2lNhHeeR7ljN94JNfcOyq0gccSMJR38tnGeVq9FsfnMzedxK
zOGU75wsPcZKTTQbKqy07VcNMmxFvvZHhEa6do+JOHqcRthbyxb2yL2v/x3IuOaB
XzM0LpT0swkN40oaDchu+lgSw+Cw1/0FQsNLqMfhH8oE5yn9+DEDM9I/XEC1q02U
ExbANjOlowV9+UUC5giu9SbnD55adIKNIDxuDvrXOqqIOqWghJhKG5PSTRCLJ+Jc
jQopzv9ivUl6M5n1CUCb1/mtA2RlqJAaq8Db3IKunq6dO5V13Oou3jSw07QVAsIh
Q376iOYKDttRTdVPCKkVfmQFAuJPJS4PzEYRgZO8r0TFF8d2FyWRTT/OcctBb1g9
yGiK+QkpITpMwGmtwhGEA63XhEU6rXrG2w8FyBAc2e/mf2RD2N8oJ9fG7baRhSPk
A2BNYcULPNwGqfT131P1kGRyJBl/24se8RRPal8p22Lcikk4BDWHEXpZXuCVXR56
mLDdYTInLAha3+SAmkZhZYAgMajX3MQI6f2xZlpikN4PuUXEe0DJWZVNfx9oAx6O
FS3hMukJNKmKRHDL0ZtiWrpn7bIYmkXniBCLX+lwgtm1HXve7j9A+aiajuPaIIkx
2I/4v1KtJIUClVmeG9IAOgJLKtVPF4qX2NPi7P14aDwhazWIXlm1zvDMbO5azou9
PgE4NsDL/sOBv7X/LN57qAXDNOMisE/IsfxdTDc+YxEawBJL3FP8eDy6LVl6gOGK
PNsCTwHcOi2i3xZbZCbWZ3GqpZDoScoBZMP63mz9cR/i0zl5Fxl3DEPxkB/ITPzR
uXefApsRw9CvGqrrzei8uGw9qzxvfpvlFUh6f56fmAvOCLN3vlV32NNFDCLClS0j
mBaIXebr2lnCdqB882x8LAL1/8ypIXpt9w4xQeD3eeqaSkaWe908/sbfr4t+lNVP
YNn1ApIPps7qM6YVt05ifeaEQAiSne3+pL3u/TZlGMPWgFMNHkEbzcmk73yqzmYO
QOkIu2jUpyrT0IxTqSiih0B3sSP6FPnk2lB9q7Xjscvhrhbg9BXuBOhdyW+BkOJw
rzQM68herGZ6JO6WhdJN09FUQEwPOhO3g8WoYFEA90Zt+LNF+9MXfhkWw04bkks1
1V3zP5qhulniVX57LcVJT5lbGj9XzLEMWuKYOvqlNauwkQBUUmXgRweAYgc1jiKu
rejAhcIGTxr8DAyQcgXq2gynV4aKb3EAekHi7UfkDMenOZBb2SHcJ3rVsn4ZVV0B
2wCJmywituS0KvlScXx4AMu88GtKdQq0YMKLuW9iwzSOaSzIb60QLCpzn0IeWkgG
3I1G7H612nY8zWOJ3XSukLwjB7Bjr/AJpDnqM4vFZHZFAeIaAWEoDmLjvKQMkgCq
cq8vjjfdNZkWRv9POAs9eEr6NciQlLi8si+Jsf9CQjtUOXSaV2sG4FPNW2Wnfv3c
Z3KF4CBudjawaNhYF4TF7a/E2OFRI/h6YL6beQuydZQGGl/dIzTZ9Li8Xod6j76C
s6FEuj3hLfdLwN2Zhhpg0zVJvZX0Da1JMEMUl/uy2E6ghk4kTDRodLZAw9u5XWNt
Uh6mQ6G2Et2eh2zpJCuxUBYX3IQ7BzMSRlLtqanfeOZVgw5AcqUbxB363aPhzTaz
kE2bq1ExIFKnNszLyTgUBTD8m9SS8gf7yV6CHgMJlrlGxy7MidteqdmiLa2EJEel
IbfR4yGuo37kyzas1InlM8yvhD+TxGDuUCpjE//L8FXanrPgPlEMoXq39I/MiMc4
nWKXfSlTRPyzgJz0gKxAcEna7+BvHhlJCraJkcXa5TwAP8k/CkHGBQZs00/4sdmJ
q9EYAJYqB2J/odv08xMG8ZlvvmLAaIifGZENKUyv8Q3HDOfvIa1wMFhtcG1w6cAt
ZwFWY/zg1Oosh0twtQKaFSWksg42PJqtVSCk0tsZjwCJ7Oq+SdJhLb/Bzq77ntte
3ne+a0tyVUGs1iOjDycEt1IZd7rNQO87Ho50amQNUTwilHeVfVSZYtmAE3Hid2Pn
eBb0nwM1IkaBQzj2dnYocFP4xSP4z9dEgEzR2268O573eo+b9PtaPSeaDwbdhdU2
vTnRkBY8usL8msW7BFhE4f0rIdCO1+mQDQnLsbVbp7jIcu5uoyAljEWhQ3YkqktT
jXTY7AXCM/065D75+MmdjNuJ5+X4bmeF0XvBEaLY0lLNzHbuMRjtKIQH+JDiILlJ
+Q9YuM4y1uVJmIbKI8Ga8gLYTyZJyBfYfghfCvdHX4I3CYP3mJGr4MFhLGWny4tY
jdzyRqBQNI+AqGLwr9an5EiM7c+zn5++ywP5L3R0NzE90ifhIvoUL2upSOngWJAB
rPIs7tDIcMMz0dMbVbt8M1iuNMBPXTF/4XQmGE9Z2CNDdaxmKwgan3gegcyEUKGx
7uUXp0me9/zC5oitp8ZjkQuAUtKZ+p95dx9sUHrvKaZHVkiM1L4FOHGoKd0CpBOo
mPfXO7X01syJnZ+ecXhwdb0dVLl5ifu9TRPwx8ocBUpAXcEdJ9SZpB8tc31ZdR9z
yI3uHQIOf0iEImMOrKp8AwYBAHVA+lcpzNjdtPGGtP9R8hkc8b1sAiZ3gFb+2cbq
dt7l966t0cBwrwhNfxxEOC7gFcbPIf9cy35NYAD5o/LQ74YkAQYo2D7acbuDfbnK
mt++nBLsApW964hlOSobqQo3kTdHhSkoij0Zh8MD+duXAHY4RiULnSVtLTYwt1IA
wTJE5LPpuBTy97MCaqMIsOC86/vLrxeEZ1ZScm+QS5dWOR9lbyZaaUumxD014bvj
ko/wWlnVLJPOlMzpJP7RE/888/OC+AuAEDXXnqk4JcnxMK6cPe8P0eGqAD1sFCRZ
lxbPYIhzVZ3VyEB1wuwrvgNmnDE/G6MylHu5LvDUHTbPpYfJw2ENFlNNonji+tOH
F98BHiJKjbSVOOIKrB/my3gGCak9w5Y/LC3FFBJ9ypkx1592mfb2g3TvTwEiOXzA
buiWxPZl9gVjxr0Dt9v7kSzB5+nou5Ttw/kGlxJ4g/JzHb4zH6dw9a5BENaANy6r
OxDxRJWemFHNFQgVt2uCgcIEDMfcRZy7PIl954QZBKlQX40URBdXpKkTvnxkvTNI
fvobvc4mjlYOSj0ozyQNEzAPFYQJ8vthpQVEMAU1s8zDXHV6s/OAK1hvIoGbEX5l
O/N9lJyKltI219eA1XQcqzctcEn/9KAQXcZ0Ie1Ud1lu9+ZfhOT0iWV7vw/RzY6q
1KxsKVlDELpbmXfBIIzfIA0YbSYeECfprCHLKRWh71Nndu4wZ9uMgKTxaNJrI5to
Vov5pud+MHuWME2gXPsGX6r7tdUTG31xUxyu0XfVr1lBqjC+27mPZT7gZGZDgWIw
BjGPcyDqxZUW4oC1W6dc5S0zzraHsEVSsOHsUIDLWtWvD2NPEspSBzKHsLIoXNq0
kWe0X5wlmwGmsXzQ0xYo1eCAMQ9j0s3px3m26tBiInsYi7Om+T/BbjwsXMfJNcwP
z0OApm6eoFuOfSXzEthi0ueajqht1+aNt087o38a1QIxLOR2lTNeHg000nK+/RAN
dCPHHxj+QKGNwNie6///2RR/Od7ulFmrdkuYluDBaqlFb5PvTpEK+Rit2LuaGzaA
xG/4b3p5ZE7vKR33Zod7kb0JlJw25U1GK6wgMefuO2xE27bPvnLqgdKbbqdxmC8z
hXpr6eDiOP+CiPuaKGm5ohFvLDSDa/fNJwv1SvnwK+kmhvytzh7mXOd/mqL/Gquz
7cg8D777xzs4rUe7rJTx55VkOrzJdYhZLdH+VcozK+ytIascD92JWt6dH3j74IVr
4eSYwgsHfYkxKyNW6KZ/hTuf4sszH5m4UCP3cf7BgWG6yKi4vv8Q9kjIugggvkGR
WOSJ5Wj23qv4bGNDtizgHt6GkL/taE2xGZl5SrteC4SvWt2CnQ4oOR1rHg8tTq2P
E741HzGxErozvtnPhMsGQDMFL5AVYkLL4QhbbHx+/SSnvI9k+CbTduzsR6/yOM9U
8ZqX7kpgFm9uRbdq8JPqyOXdFIZadCXuTIqqRxYJR/3X+R8TD2rFP38O2H6BgHBL
78Uw5snts/wpZXiTCzPTaEv7Tjjw1GlcVlf5SeKu64Wf3C/nRRMoHZHcVvv7Ofs4
ZnuFFNQMcyjlVPApMlgk1ZiEPKwuVwI7e+MqqwyJGxttJCCHa2837LJAES+vfexM
0RkJ6tIlfjY3JoCR/Yhp9VK2NbD9oaYt0telC/9g8GOjMf203A32030dzgm8gi1F
jpuJ1IFhmeB9hge/bdUIzWqgBQOOKnZzAlumtw/C6+7N3tTlMX8LCN1SdiDVwT4n
axtpVzqKGL08iNefme6MY8HgZ/01M8AvBFpNcaYVnOqB1lZhrH5w8H8YBe6ccGSt
3/u+vKOFq7o0sQmvAdGLfu75GmuRC/i3+oibSGMNjg9QyfKc5qQ2oYX2HjU9vsGZ
J5l/uZv28czg2xiFYbtw1wm27kJaTWFg2tkNq3gfjAyZLIMkl614z/Pw99Mzxi+E
M3jRDI8Oger4ue0ejlnRQyet2CpTgiozJDzY5aHoaHJ9ImOINw9e4XVdEI2IdZIy
4RW3Q9OuRdotZrYwdF7qOWZqAKVBOg807tCa0y4VGBHUA+0njeHbPm5srXp26HoG
ljq0hPpPCWaj1P9KL1GUfdKbeBgdSXbQtaa7NesUc/+NAd4t5411MTQK3nOR4P0K
KWFQGTQeIZ7ddu5k4Y6OLWhQqpaK5mmGOf52SsTRM0FGpd7IyoFRnoS2GlsJAWG5
4wdZOd9EmyIICInYzYBaaB1LoeuudP/mWGJVOpqmeL36RkgJbQYlr171xp2GIwnt
MfLLoDLoMCoupULnrNuoEWiGYoSE8PF4ItXsc/atj1wkUwHjsHZkndTsV33ii4f0
129wWQuiDdXdLp64gs5fUTFrOkow8SaRxL2CRJk+V3Gp8+xHAK41rrsGu2DbuouM
tcP8zYKSgxgCp5niK1IFdyAdZMqX82TKy7Aa19kyXHXE04w+V8C4iUwuI2fw5V8u
BxnpMh9rJFvvJdjGpbZH6aiKah0hKdqTZ9P7sU7ZwRpXVQl1Q6SutnByDvUJHGPS
UZZ2U8SHIlfzCa+Sxzy+LTxt6VZVtOTHVOI6p9iJt0bf05mrLWIjjhFlbMiRNVFc
jfHYbkTqat3vsi0sZpt2MKrv0tUbh/x40mmBxs29jwQj3TSUPaBpHz/LigwYSuC1
Ri1FBvPtmhqMjCQJyJ/BEZycwYQWBFzy7JWzJV1sYyh+CZt1MUZItj7TvsnFxvuw
3NkTTN/GF0rrq+Vqq2/f0sWWajhhAtZY5VesqBbwWL/DSAltsDBsyXI/oW5QSr+o
wxS84L/gbX2z969Jj0o+N8Nu5rEfIgPhGYyqRR1gRlqyQxesbaw+kb9DQIl7sKxm
QgADOH1OXBBP56Lx1sXnDk2FrvXnNGdkzPCscTWrQOIyxoRxHaIpGSUbZkonNWrr
tXGAU3Pfx3PPTH2j1XHvO9kcRYmHKHJeqhu2syXhbHY3nHUrQ/lhRfOPlCgoKWzt
xlwQGG0OEGWg4HZ4g3sQKln9yepeHeH+EDq0JTF46PYSBLMsH7CSUksoTYzLqcdT
9o0vs6E9TGqsOf1zfP67LmYWhspGhYPRR3hNZn0innNsw8AtNlVDELw/8TODeURi
ek2qsR51Ny0MyHtS/qEY7OB3sTbyRin4CfzQQuvBKbtSauBbsZ6IvywIRUZAbYaD
6lbTKXnEH0QMFGyHOAopY75SdI6meESUF0XMUigSwwKdEZkc+W1yNrYf13cr7zam
Zw+e+jkia4/00OtrdID27T73pD4psVR/h6nz8pH6mnqXNKhKH9NGgNc2Vbwqt0/Y
w14T8MBX/TV6/uEB0mJX2wLC43WmVuWr0rLdQ7e01I82HxxDgZbFsKoVfNzb2SoD
R13z1yNpUIXY6daTXipKg68jiKs7hE2qtAjemdFpEwfD3IRwdGWDuXN8xyceCSxq
vh6ojT65ZcFZnv0RR58nTGCK486XuBWTA7RjkvcLgiK55DdvuXMBweLBCZvxdQau
vii57PGUwOuuVh0TJPeD8U7l9zzH+Yc78OM77JMsOfW0puXZNoZfeGlomPckua58
8U3kmpwDKfUuRtE1irSbv+T8BwFUyouWuVfjMXcemqQvsYvepSNskTD7XOoBDX2K
8HPKY3N0JemPdXVlRK3wrMxpwoAVUsEQfYpEjmYAtzzXsApx8CDRs4Ch/oewpi/d
3KrLa8fhEqu+8YIP5nT1EIUKWNJcab3caM4KGQsz0yTTaRElHFTll4ym+FvYtIfW
0cRSLgcZcTaytb75b7IsaVGd5kr7tDaB5rfoV0TMlerqcKlTghS6S/mWj+NDiUxN
GnUwUvh2a4BCIQ5O0CUE1WmqgFan+hxOW2qE5tRVBdwEvYB8AOOquoVEKMKUDpJa
rLnvUMzifbW9s1n70shMrMUX7oEJ5fhYkgH+1uVI79IOxBbirRhqadL1D9i5P1H0
qO7olFZJ7MxoBwDrudQFYN+krF81KyeaXuf1L2rAUw21vgE+xzYPYH7wXxNUeVus
A0TDVx3ED4Kt/4WSXDOIIWzD1OY9gPQ0zk9aH+AvMHXqM8s64qB9YfSfReqA4abS
SahgRLJa28IzPxtr3kWdYPxfFKsHSBibXD8yxUpEboq5TWUoBX83Zb+WYV5Z3nhB
4VH0M42tGVBBj9BuoPBGtIprQGT8ga3VwuJlGRSiZGiQOgfyYS9nLeIclMphxdY6
PjwmIUpxHIw1W78NR9heyy2D4Xyi3mDR9NqcfDtgMe5OJWViPHyeyobU4xx6B/fl
+weQY91wUGSGXX00Zx90WHri+dwadOe+wzXR5B4fSsbR6xYIbyZefqdTFBBy2u3X
rgkt55hL61v70Dp+W6ztEBZCbNZQlV5pENY/5fDwFyjccyo0rWyrJtNG9ScQJCcB
GtY7E3ucK0HnpSDvpz5tDgEDFBxy+mVX7a/eE3aOZUaJ6/KTFjASGJVZ7Ow5aSgM
AS82+MhcNakcYTWMnkRKu0P5E/dK0xW08B3gEXYEKlaGO/KLsQh90i+jyVGNnxdO
LGwdmgGXMugBLzk9/7JXMQEuRvFQwxkyxtqBVnfT00pyROkyyO34cDi98Vc+m2Yl
agn8XtOxn0Hv8ZZP38vbWDEMn0Cv7SmdWakCTMIgrgBPRhan+wPDLrOgHTxeMMiF
oSN6Fc9GUbxkZJAPWPmWdvG+USohDvDo0Y/dqBtbk6dnz6k+rG+kfSwLfLKBcGEM
ss70DxJEANiIN5kQpHIObS2R5Ps+vQIS9eL2zCjqgVcd6JzSfzPpkdtl4gKnEkfE
RK6JQM1yZjv21RTRI/pLbCacS1BR0k0FbKYjVWAoddX4OtoWj/VLEupfiZcLWMEj
hzkUU6XY73MZCjSf6ywgFlhrfY7dY3waymWAxF5o8RSjKRHz7FxvGuCC4VER5biQ
6GbEsm8YjpfTfDIXnNoIlmlhK5+ADX1UXeEIpw0+Th1j74q+nIhyGmOHYFtFwqnJ
Aj5Na3KqWFIraHQtytKTgqPT49rQSKDv/viDpfXY0u3HbuMSUDTfgQBCQAKDEYDL
PO3v4muYBLxF235FduENNv4fe8vM8UXFpxTzW/LBRetYxOjN9j2pBSDnKW9MjoPx
3/MnBKZyVCzGuj8e3iQrUf0qkCFHFwCUmZZlCoKj/hm/8cIyArskJtR0ko1UvrWV
DNvowoADHCWks4loyp/ztsFZurN/k+sfTIuAa2t6I8AYV5cykG8vQ+ZrRPhb1Xhk
M9LZzWg/a/N1ERKkkf3whTFlbzTbeSxiFuK5mBM6cd/k0BCdYdKMTJmNzZiQNCtF
aeNHFhaJGmwFLH+khvrEC6lHRynB4D5PUXi1nP9F2gy8fM7bQywn5KruGXIZCcXQ
YnBj3qqypzWeS41TI9Mmqr+cW4H7vGM/PB4VCwVJBw2RmHZLxR9ssPOVklPFgU9U
0QHpzODJjXzoYaWa/gnnNshpc0bk50MmQVAsh6pzTG6qb3Abrng+uxev0S/LnbvW
27ct2/F2ogLpk60aYTPGUxybdYCFl96TlZitL01PTnIMICUj8WSApG+mvgQev9xj
W6jNivSrNOSm6M2RcFIX5C6gPyIyRC2hcVZEKv2Z02rKbqQfgwauobESsRadtlbN
A/jzBMQ4F7i6QU7HQDNJ+ROfNnNJD/Exizxe5jRJUO00bBDwldcXAzIciq1ght9J
WpwaYGtjgV+4qUw0DQM67FnlixB36u0N5dlQw0ZXc1z1GZlipQgFjofp8T0ZGE6c
USoqT+nvJnTowBO3UG2WNeSWok7JNHE1t9YlMaJU8tPLDy3wtWZqFG+/xlgRMXzV
cXNvwYzWIAhXujBzNNccwHQapnQB7I0ytVm+qy853U7o+lanLBujguT+3Qvc2PjA
0S+RApPMFqsucJCW2G23fh0ST47UZYzwooLN364RlE6wUs4pA2yzXsd6fDMBWO6c
Z4H4KcmMQFej8AkoM8lCFB6IwFF/JRMM1L7muqmfGhlldl/1JOfytlNs5S7N2HQn
dGVVBXn7p4peSqTC6/8HwK7oOsrNlOzmXcjaFXPzsu7XW/Aafx9T/OWt0VlqP41Y
tdZmVzUWHpED2KR366HcFF5ywVskQ0Cy6ev60kO70lgbtKRmI0PUXrKof8FtZuul
+/ozOKZgCqrLuKp7Ycc4KZVNJ632xhaskHPhSUMcAV3pa8wwJjbdzIEldHNz5/KK
RyAod7QtdHiUppxgNjY47P4XxTJujSOLvZ6MW3FjuB01awBt0Nk6FEeVvC6+05xG
Ar2D0zUl4JS1ceQ7kctoeTcuouoDgKo1G6z6AG2iZDZI4vyV+uS4E6SUlXLNq4p+
pvgHeQmo9iVW1SJZC6ayktJtOd5PX8p37eVF9uxoc2/XT++LQErAHEM+mZT2lrQa
fVKcC/gYMLreGsm9DKF50c4fAxWjErpqjQ0etaX3GVRg7GBHVKXyPKnNJNw2I1Gu
yz2A54jW06KTVcGDM1MHN82kJRa4pQ640BibPsDRyaZNnbjRksTSXfQ5jpIAxw4M
b+lL4x4vZkchTn0kdA2jZtezHhsfXLB5BiaUJXB2US8cW2XgTw6cOcbY3AMGLAEP
mfHZ27bVXWBNL5+4JAjmFuziMsHNe+sLqmPfnr42VhLCg6GTCRfydPJ7Q+Ao50Sj
VOd9NyOYKmHYrLPTL/nN43y+JjdcQPGSfWu8MhdEfYzb+iay2vrluMycs3bEcHNQ
H2Va8TUjlQbo3bPF5xoBW2d4YimBjJfes80jg0Z4le20CbtHShwRnkpho3J2dLac
gd4bXqUkYhg17AFaXtgfCeVrGMGYQ9Nhgr0sJMKnN8erjIW8TZjIFrqtegxtwEN9
Xr/AjtFRxcsMVZCpNsuuYIuia42WdSKzQMKBAloEszmSjcnBGJDI0IpG+S/eiw6E
wTmrgTLQ+tNxh4DSXxKwWYNGqOoM62jrud+R6NcdD2MKjH84esnssQg/KnLlepid
cxOUOo8JBoTQPR0A5ISu2X6Gr/4/H/yRdi6VLTwZx062b9AO/3CZAYNiwH7cSbSs
O/GSkGAHP1YyHEhx2csK4k9C7RCOXjKQYC6hFJeFBVnfq6Tx/4FgsD4kzktTLrUb
K+8tba/rz9D2cnn0bnyWlQ781Ia5MjTysZzulBr+FjFEdlZOOg5udn4V1lZy9xzn
rAVp4KF5wJuu5lJE1VV/W1vNUNcsEzWYTlXwMkvM8KYq7g19+eCK7NkGCl4VTve/
EJ2GUN8uqv+pI7XmI1Pcis0doAfL0qd/QAbqOI8KYVRGAZvH6kAr785pyfO+5ioD
WXugUq60P1B+HXjrLSg2gVB9ZzTVmjdi7vgflZ6Fsz4EV8/Vke7nTM3TcW6V/QB3
/PDs0dpzE3HxSl+sZqQWwDwN8SA1YSGvvewYM37/N+nHiGZMpiq8DURKLTzWP3ar
dizhzoMbNJ850+GRIfZ7NM8fat1RpggiaKuxBVzyXMkeaAvruxY0IflPk3lgvJL4
byKdner5nFRO3lkpLKIxgc/Su35/ryOUBkJvTeYGpO78DB8QKT/xtnAVSiBFfiKk
4GUpry3PA/K1zShQfGDkqm7Hxg70fMsMzq7qr+Hlw1ZzW4do1UZ7y/8a11+97aeH
frxHVH7jHxrWosY9zebd+0SUJjU1d0jLhsTAdnu4b2RzBlMzMXdRsq0eVMHqnJOJ
aVi3Z8V/l0IkqOOfLljDqcQtbdC6JntzqykekF4H0pIXxnq6lI3zuC6xjmUMDAMp
J2GeJpkOWYh0YEmOB67CZKIECmjAEWbD2DsgaLOFC9oUA7ZdiGSXmTo5PFVC2F5u
4sQwb4StKw4NKW1P+2XggoVovnY+gCdfy7yvZoKB/tJICXj8dYEiehmHeSJZYjBH
wUR4Lz7py0rClZeY9LK5ZPAJkKCbB7ys6iqLT6OH0IuJg1v7hIlBjXF0q1vnzrOS
p0zJJ55OYYXw6Gb3XljT0UyJBT2n/Ev1+eBU8M1PBQs5u/3ChwujpPvB/19qwkd4
sr7Du3RQvnSWJukPBZslw2CniovV4MtHDYckWINY+ggJmdhdRXTIaGWgCkiX+lg8
yfW829EdnI8/htccwan8oZadkJk+5MsbguJUq8ZX2r5G5Y1PoeYhCV/eD+4/OjXc
IJrb5b3ixDZw8cJ9wLDjXFU+RBqny2zoV+bQLjPSpOS2ilVoQBFGpafHrmQk+coD
aXzSNny9dRs46qEzoZ35IGjYslRIyy09loo47scDDA+7nuuNT2KJ5vpM2SzRn+1o
Q75ZUSRabcAHLa3TP06nXDMHOiImoXvdemozod9GQOAqCWcV1RleOhikjRPMqTOf
+0Z+9U8TSCKfZFLE4Lu3H/kYxsxOdVRvWZ1wU5lGrhUR9Oaa1xtiIWWjCALGUplz
DBtV5qsERvD/3NzeKGzqA0PfM6JO0Yp8X7j+mjq5mKLVg1KVQ2evfbYsZdhUk9wT
8Cix80ZwcFsHC5qxEKlIW08K4XuqNDL+1IJpx9Io9aJG6J2f4fZQTl90obs+VqIB
pqZWo8FfQfGsN6rbX1ug/ugnMF52RB1Rlwh/Ayw/4kQb8eAK4M1xreNRIIqc5dVz
u7R2bOnpp+DfFcBDd+Yox37yfzHqfp8KtLjxYBHD9F1Tjug3s+7Wp494BV7MS1Te
sJ9t4yOuliKuJXGBtYm+fkUH5sIFQsbGBq01G6hK1YQT8wTOQnjSJSjXerltdJHg
h6xsJEJo7MOCxr5RR2clXIjg6o8AXajsy8AKMOMV9nKeWsjpUqKDNfyBScOipn2F
TKvQ9BGqt28wU2Ok+gP2eM457Sg+UFZhgjvyAgkOvQFIsqLhfbBe1hHeLbeUgEQH
rBT/lBsIYQlXUi/RsT/w+E1rVwD7uMF1TBkXXgi7l23OIHkQ3pcYgLRJ5/W03sLk
9AIB9wWY8lfL0EJUknXXokP5I30pEn4kZ0er/D+WVAbCr8Ji0pPunvkARr/RJzsc
nbg447LBShos2QEQ9XddrHWvKO3ejL3ZADeOrWscHh2rdxXHZwPQBYXIE3F9ks4i
LgLhO/TqkN19sTSRTqp0n+hh24/IGNIaE+ApUMVHKD7NSoDE9dZU0LqDW+Br4fz/
r2BanxXjZiv3FwFASDdz0R9q3xJpdOQ1HBNqlThrBwnYXsSnEQXL8JlAjuhn6WdL
GshE012nlmMqr/o+30RWNAVUAI42vj8RwvaG0jRBHixJez8o8ralwFTRfcr5Ilj6
4wp/Xtp0FbNPPbJrZdmn16Lz47PIJ61IgLPgphcoEtWsZUyu+FYzQmpWyfmJzrRe
akuVp1XxAq5xK0ie19NL3t8CC2f+PfgC1kkGoWvnLBTbcrNr+JJiUksxoXRQfszG
nswoaU6omrUNC1ztdAfpZAnacvavyad8WQFG4lILn9tC4a1EIPVp6o/A5av0GYsD
xNPlDJ72CjiheZba/vmQXZCYqKaABsSe0un++vL2WknoO42IdnMNN9zfU+gtcr2d
7qbNbtN3GX+mckhrK9XnPxYg7XCJj4l9de4EZagSQYXuXSRO5LWBKniDcc3KcS34
qLJPfx/LNxoZ41YB6VN5uvOAYDUkR/wWfchdIY1M5IM31J+GK3b4btZpknKXxugA
zVYQd4yT4YWOK0JS9KKFtExIhvj3qNWBDkF62wlTvevUNidR56CS2qXhPlXRyMDx
WRDDxVnvEn/C6SwLTAdCYDB85wEtfQ6HL8/6FgP6YSArg+jMGsWWfbzDgPR9NKQW
7w3CVSv9V0J++yHRdIvYVP/2UJ3JWCXIQ3RJe9sqdmj52ipt2NfOovxOMiPDNR9o
r7TlmKAL9XH6RSIvU6uFuN6MQztihUbcvqqdOHKHNpG72jTWHQRtWZUH3BdRQKcg
KJgJFrV/vdtd0YgXBAd/iAj0dU+n5TX+Z1DJhg68+VDkYIzywPuN7sy+0OyivTvK
3HRrxUUNJcEyU5aIyPEzo+1sWRA0WYQXSdS8B4wZOcqiBDDBSVlTjMq2O9pGBcLR
roU1YrJLikbYdgPE5eR3SQvggqq6m/AOg52enjNTuayGijph7l0XxHtMXDNRNzH9
bMYe/WyU0/UXAJTxoHmqI9MVWlY0bjmfrSuEraulIgfXtLKa7c7jHwYLNIZfuJ3+
x0e0V+m/c5OmE0liWhPhCrNSVOy7KhlS8Hw2CNniV0YbxzBWXcAkH5tdM+/Vz6dY
UPs67TZFN52JHGKgZCcO1HHT7KoiKSWpfw14qml8vPODfCiURrkCZnh8Up3OicKG
7pScBKONws+8TFr2/za+cFkj4lmlIrmtliGqEfcL6IdEXHSRwgpnPWil4l/SQgU9
lCfC+bMQSiWNi1QUAdghV3HVUNQbZsk53liBcY7CxiiaWjaa+zNgKIWnHBCxwuDl
V04v2C1H3ooG5XcA51ayUhI9+HauTN4inuXREie2KFVSr4J6urz1DMUxUZUZ9sm8
BPLGyDnZHk3yo4Oc6LQoL+h97caldG3+dUeuedBh9siO8BqHJvCdcFJveloC/BkZ
IwjcljkmBbNglJromWlddgBta14enFCseEuOK4QYwA9KubzIZplNeGdE05WaMjCk
VcZFQPl3s3XeddsSzbUkTWpI6IElNZK7knjXKpwUmHLHaK5y5i4QDegquaGCreLK
hFtH/WO0dzacLrs0BWRCpaWmImR20+KouBsYxaMKbxxRu03z1vCmvEsThm2m66nI
6L3gQOXlBo+MYlA8qnMzG89PBh5yeA6vtXyeOozRVP8F01gaiIx5ATFOdzvwmtaC
gwMqfKcq0Yl+yaf002bRswgOgcAA+sJ6rbFO/vb2ayxEjW7Md+PqfwiUTQn8FRbP
C4DOQL0qNcIVR+fJR9JC4cXVwGUTS3tvBrR2FFDkdDAo9z+TJ7fpk6G6Wh4bBcbS
gseLF+349sgcxCjkuvUzcYHNY0EtAc6a5iVheF15H8/Iz1CRn9YPNKOb4SizMkJy
s9rGgknSVVAQeehz5QefhjeLJeDLENjmLWXHCUt6u/3b1K85UOv9p4pLLBaWiJ0B
NWQXTS/hXTZlfjrdugPbzZBIPqL4mvctZPT65PnIVk5ANoLKMlzfNdYMtTMAw0Cg
Hy0+2F1S+mTvCqoNvI1Ur+MAGPG7TbznIRbncikVHRoj79fJIxNdgzzCpNffDRWi
dEo+9KVI5ynXqRQE6WcSKZOg2Z/pL97zZ72pqjxzH78IwPL0HmHVnigfTyjegS2V
E7qBuk6UGaJFfnvlWqfktHEWCHf/Pf4009dMZ2jZh+4MHS3bqkV/DLPPD5n0bvLk
Fv8Gu4Bq5Et+gbLvAJCTkS2eUrW3cdV2Q9cMVzXB27i/Pca6xqims9X1Q6+zFaU8
XUwY8oEk44nZd+0x9vbI9Veds+NDXMqut/yffapaOUp5+KNMgpA86oQOE4OECbr+
WFIs/1HCnyXsPtBT4LF+CBRlQprf5v/l9dgthsa85KXihfUQs9U+ed75WKIWjvOM
z5RBKAOnrPUNu6WpeeKdghcew8+HDQe8F7YadzsVwAxmmw3k2QkRxGEHz7SNu+nf
bHDAwd9V8gsvtXU75wKFxpIcajfLY+0aZjf7dLTa/zvHNOWcuHLeAWl5vRXkfgzj
CrMtPeFOba/CBDcZHcMFsj/uaDrafKoNVsYq5SMpilvOOUBSbQT3ffssX7yKjbW/
Iqme1vOL757N77ZD/OoTONUXCPZre7UEE/Daq1eVSAHikbWGVQlFBReoQxCNY5PV
BRYVn3SVftROKY2Tc62hLV54u7OhvTqBuS/GiLWTl0/TaJ5RCrCemFRlTKGFw5ga
0aZvEym7v/htawGVZrKUNgS4I4/lGjMrWe1X12350pbSaA6rdPMKRhYd4DmMF4Ox
jw281OpL2xZv0Af9T3TchUdCn3nq8zeZ3Oc0zWT0C9BB4LNflBo1zekRk2qEVF02
SxYk3c5czdHQDgx9yNuqj9lrhFebiHGsfpziDe70N2LyHe7TSNXMYqnEzH85xGRL
f0ueLeDBTVw6IvVEq+R6mQY4yhRM21buuRl+6ikV1bbCJ0ZHryrwSqR1X3DQjT2i
lyxHQ5wzMSu/qwyOWSUzB0aD0hrB4fZLP1XOaXk6d5ME9lgvgeNJTIbpMSbQAP+g
iYBPTHUaX+HLSzYriNf5XJVdZsY3zhkRQfEvXSviTN6rBm5LJEGn2VxoJaioziMz
QkEtCHkefsln/6pnzdHZ5mCsba1xo1DJTOj3jrQCTC1HI/PX/Q9MYND6HXVxDnmK
onntCHJxSu/dYORE79pV6WHvGQSruRXtd3s8DoG2cAmc3kXmOzgHiLeqUwsYdXxE
EOyX5NK1RskhEfPeOOQbmLBJgD/L8jKhRe4yx9ECkUlhKUBSzkUwDdE33lycxsA3
gmeqYTlVcxYCQJmGJ80m+QWOVdPbBInDs7fyC+tlB2ewWJNjouM2enkqHC6brBQn
Y3GwiHepDkySp+XgG+TGUfTmHJ6gbQokD9zP23MlfinnkxefsPBCM+k2nOa3gXHH
lcaPseDkEm2jlMoCX0Dz6pceq9KZoh9uH7KPVN2gbsribdVi9mA4LLqgGlA27wYQ
4wbgk8gOTwOlGEg7JipMTOcX14ZoL7+UWlrkUHe//+rQo/ubeHwgCXORyTt2fSbY
oBiUJaymwyHTAtRVQoxe3rwnI4/kODFYT1LVrfb2c8QZ6xEMstjM9l5VRtZU82QA
HQL0FxNplU2DcS0qSlDKmvbPWpzbUCeIGdxu2oRgWEit+bOMzUWHGhzHa6TpmjAr
Zt0xZtlxjtifdQ+0zulgPocnJUPXtje93nsaWF+UX6OBErCwmLclvCyqpPg+4K1A
2536DoG0Qv7LKCU3QEA2JG1Mdv4YB2PzxIB2RqufhV4=
`pragma protect end_protected
