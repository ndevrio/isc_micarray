-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
G7JqARgdg2XmcoGxB6pq//nX5FT9vZpsIKuKrI+CtFJ5JL0OoV5qa1UPymh2P34M
HrF4WPCVGjUSEquk51aAcFlk1OOhRLAdyv3TWZJlGcpjYS6UZG01OWg/Eg8q8RmY
Y8eiZqyUQcfVv9DcKWAYdfqEpYV+ZbYtPct6xNCz748=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 2549)

`protect DATA_BLOCK
Ze4JlHAKamOovbljv0sN9YxHAfFDSyjwYpvJ6MkluovjJrbapwjfcrDPweCFPkbq
yGJ1CyAgUOAVKbK/GGsAa2OjS3+sLwu9bolcdmOEslZKT1m0ktA9pPr3WwVbePxJ
Ev4gPvtUDl2rxApTrI4ka+AV9HplOkhmy3A78iIXH8ItrTv42fuimnnovdWh0CvC
x1PcVhYywI3PmJ/7USX3X5A/mlhImL7Ipu9e0Wrkh81LTA0uCYE4pOf1PPBclqyw
c9kyI2RXcMQ69opyVd0k2dXREJXj34YKmyuQZiK6fah+IfplM+fVWR33ElCcuZ5e
kQ+4x1MaF1BdZMcdSI8BcGLUpM0qIFQ/HYJNOmitey3GBzcoeKqKC439mZgreVhZ
BNQMm1BIFlW9AyrGy1f/oEtSR2K3GAuloXMzRWOK7KZsWIDQNRRGYfA25QoAB5Tq
2iR3NsYGo2jCUEty+bKsAtcPFPUG4zjyrxf1KCzHv+lSAtIcuQiz/+XLRUYe/ccV
tWPBsp11Q0oVezG1skmod306+PjZ6WZoQTroREewIgFETvZ07QUgsqHSWxSfsBTi
hCN5O5H30Dscwk/nOXw/aGTpQvggMvJCX2M9AjKqGxFHdEkwjcWtVX6Su+3Aq6GW
LPO2PpQSZZ0NGrv8sG0UyfLwxVZ5Ge5anvh+5qad145gPgsZwosrEWdbddyVA0s3
pbIaUBMn9OkT83weQOGhPRJpSdv+6eDUeUU4h1WMfmkdlMaBzhkH6eJ5x9Yi4ocr
hImB6A1+j9fBCkrjMbbzgAx7yLbO+lsw3EML1TD8SYF9dG31jvL347YyCEqo9AcK
4y4i+f2VgUNF0bw2+oM+e+OI5nF6FK6X+K9kybuumItMDLNpSE3tV4CRfMFssO4O
m1za0P3trFmdt3Q8jFM189XF9md2kqrc7i712rrvD/mugR3W+X9IHyKhvU4HW8Sj
ZBpBrWWB9leSuvF5qGpsC4YkNqxf8KKeGBn5eJc5XTlSJoqyQ0KwN3RBooPQ0Ves
y9a8PNVsKYFgYHLBmy7U7VRlbMmp1ql4NqWUzGkXj3/0g83xd2MhcktGrQF01Zev
q6KqlqGslzJErJdIH7sEbKuQnivgK96LNQ5wka1fb8AoC4Zc2jT038fEI1Iffah4
EG8UHTf5IwLm6oJU3bY3j727Q79r4YF5YV0BilIb/dMhbDWz9lQQ4htxY2xPhP//
MJ13mH/AfQ8py275w95WG22BlxUJv5pZ7lbPYTgYxDP++uo6s333mkTcuK+TmirW
38YJCR2o5t7h4x8oBmIPyYUA8uArgtOjQywWSifXZBVTXymSln9ZGvvVqnf0awYu
qhSaXw2SbXCrqV5wukFqDY6tNWKniEPoBUW/PR2vz82MkUhAgxG5e9Skc3NM+iJL
Hfu1SQalAZqEOLXOzXR6n5ls/wxvANPks/KGeIMdBqi7d8tM3zLhN8Fthy3lMlEU
WnFZD+WxXlvTM8rMxSmWQiB8boHvlySKKTqONGIu9IgMSQ+6c0oVgpBQs44/8ZQX
ObuCz2iNYd5679jXCmZfG2Tbp7G8SYNp5fgwi+40cEjgEgHiExn6EA6RGLSadBv0
s7ESZKpINFF1LpukwnCt1Za9Glt/HxS7AqglWKpE2eXvPxQ96XDllNELNMgahhP3
smyGKLgPysE+efAHfkUr+FVYqO048U9kVnXIyjZozmkqy3CQMuuFSKgL1Em8fTc8
6J6VcfJ+cwGd0htlJkij2Pjb/VDRRkaDmFKXr5SEBeLB0Uv+cKaKG8NGpXUj8n7C
ixkOd0g90Q89rMe2FyyaXtdJe4Iw3MXANE2+hlvCFxYXTxJFtk6PgZAcXzvG40wq
snYO8BREfxYDKzF8pIM0iKSUDHtsf7tSZbrz6p3jZDZUniV9umhLLRg2Llf6I4jb
BciEZ+WK8OMK0wYAUxj5AdD5qvdWaOI6eq3RY5lGGqUgwPMw5avMCzP/dU+sszuC
+cgbmN0+NSXebS943LD+5SVsGvL1Cb8hKg9QVJNryDDBjS9625+jROSbih8lvwv9
CxR8AxfpL21uU8LFI5Dl6dc2FS6HafEw2jWtjUJtiIkwsCJ0anj+9fpBZNdkgyuY
6UsIjzuOWyx1eVG+oczdn+Ueq5+EcDMDS2VRgvNbjnpUPP8nw6LkJNXcovk7mEN1
jnQ1hRYCJDRz4rK20RSHnTYmfUW8McPXejj7qA1o5QNUW1o75ykMV/Peo7C4JGr1
SkWAmktJK280xamVzPew8jQZtEcInD6dDKx+/AqIeGmReul1MG8cMIlfS49y4jqe
H2P6CgFg+Liy5H09ah+TSlPij+Kf1wJXx5v+zT1goF1Lg6eeC7bYx4PZ9DKI+c3H
9J35tUmeXQg34Rmlj2m+6WJI1e7AOseM1ih7wLDLNemHLh7Thvou5bvq4qe54Odk
0VzXRMs7Zjak8ehSL5djSHwcMqorFa4+qiH0wGyJdODita1gX2cE6GTEYHa1dM1R
PhORbP6TiM0wewjDIq/Nl66mBO3o2Usd/N0gA9NVmv8nhgSAw8qKcErIiJXNrRd3
UhhKqorb7c6MpOQsQZ6sEHfW/y59z4n7owwVQXZ6tVgFNw8c/FkjF/EPmeV3C1nM
OwKE7NsAKJzXQZiQLqifDcq8UTPM/vXCpW+aPcuPC76k2QhRL8gtRQpDGH/e8S39
wOFXgtPofjziww2oqEvXEHY5qTIa6hmsjNPEYuSRFrGbUunt6AfpsL4hYbuqehqh
3T4yR15zB/tjSxLWvfstW3r0pN++WcAwnHEjr0RB3WXWnWeH0cHU9Pdr+9Hpsz6H
Hlnk+OpbkUkM0yIeDxqdroHeLypPhb1Qu/vzfUiqypn53133mzR1ae0sYn4u34C3
wO/SM7EeemRyZ93kQCrY0crhH5tbvd81V4Iae8LxYsYxKUMImak8PzXmVPwnxQq7
KhjVfAXFzMUq38cDrm7AjS+FrOu11zc93pMP47klPAU2Lx76dgVZGiekBXO5vwIN
GvjH0ZKh8U/NJM2y5qnc5/BXXE/CmUsmaFWwv5mqSjf/DFWem6gmKhi9Z0+6sRoG
dqdj/XiwmtQPcdq6VDjSaqtiwzQTmnCh1UH1qrQ4jKLvnP9ZpjwBRtMCDVKSS1Ic
d/vu1rmSNuEipmXyUttT4K0GPUTfCNllu6RD5oVhJwUD/xogZmi2QjB84zpyuHIk
c9JE8c70lvlIo3jSDRGZbQGpW6n47Vehz1w/IIZnnc1jCPGrFpIImWpv0wjCVja9
jMwoXcUvqNK9imEMEypYlEZghEPiHqvfghJqiOcWu9FdiRZ7lREdwh6kR5ZWsW57
vfr7jU0dYmn3abaRmUCcIHtn8dgHmOHOQPpuyl0y2bhQ6XCfNtT0A9dEBDT72dZk
tgnQ603mqnwvFqiAy5mC9YFJl/i4g+jiIhsO53KzgkY=
`protect END_PROTECTED