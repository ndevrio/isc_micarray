// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H%8V\)T@)1YYM8.,MBGN)*TWN3BZH_D:Q/<?S'^421]<\1F'8*:RQ)P  
HQ8P?BK+9-^'CK0J Y6N5/Q\GX1\2TS^E"V-"%\33JE/Z7L/I&$,V&@  
H8%ZTS?([N'6V3#GW<5@#6$2 ?D(@H)C77*PV>>N,R71#AJ1.5CZ'BP  
H;RNR(JYWD+%U^_M*]B3,<<.&QJZ_Q,$\6(&9PY.W,=4MO_DOQV_BT   
HIN)5:+"Y@(8A3D!"(#)J,2<,V9]^7)N^^KMNSM7G@Z C J5I0*="X   
`pragma protect encoding=(enctype="uuencode",bytes=18896       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@'X$K3RM@ID6XVLFFT_Y![^W'3<I,)'FOD7 W<8=CVY, 
@ZT]--P07."12A;Y&KI/Y."@=!F[XRD,DQ+/*'<P X'D 
@+R:%)T"[PVG/4RLG^F+S,:#<!RXL^A19HG51[.VPS[  
@2O-<P!+PE?BE$ @ZU06=P><NHM^)3K?XK?8L6<_-W"  
@'GC^&*0/*X#[>PUOL5;(<1[&#ZIH"!@.FN#GOC)JSN  
@?PM<^7.^@;P#&(:L DB\$!F+.8U78A7$,$*G:_MQXPL 
@U38A8,^CR 03<O=!%#B]=I*IA7&U0T 7;/Q+Y5)]\AP 
@0.?P*G#_SQ@AE?I"[4;>0*C*OB.> <G!++V'; 7,"-@ 
@$_EYS0^2!&LF'FAXXQ2$<;FKJ+S.\TOG$C%P/N-%C90 
@C"%^5P6HO:0WIT <4.67/$:"2TCX!H%0#JA;&\:O_4D 
@V\0Z32;3S651H1B7_!ONP.I4?'JXI,VFZ99="4N4 )P 
@D/>$JL12)B-08.2;:1.JJR\>_+$7>N>Z+1=D?<: O:P 
@FRM-7'H %01)HO.5I#]^.E+3YO;S=D]J+]:VV=6"2SP 
@WQJJ/%$97J@_)A^#3HZP_6X\);1H.S_057:%GBHD%*L 
@,\I*CI7YR?L4I5T.@S2?&R9J11<"PI2=H$[58NXBW*P 
@4\?QZ1WV+S941P*E6=R<8TM-IWA-4'6<TN -M3L3U"  
@U18E-ZQ3B%B&H?E[AH6!#I$@U5*1NH+L&&E=TLI7PT0 
@CM3#GBH#I$BQ*R7HI-FDBZ,",M!0+-<X?U U9;MV1E@ 
@Q7:W[!EW,>I$T^%+FW,Z3L@E4X/CT^MH4E8DJI88LK< 
@-3DE"$0G*NE.PXVUH^]R$3+6%U5>%-BS#M^F^T:M!S  
@RU:&GV"XC.?F'U\Y>GNR<=X'27Q@ZD3\0Y'5[H>I^,4 
@W\8,Q$\]O3]FW5":M5EW(Y>B]/Y$HV+<W QP:VE3X+\ 
@2*<L2!WFTP03EN76T6NH,X%Y*K/> B"J:?35BYXY/48 
@88&1COQVB35XGWE8+,;))/ TXA"D6Z8ZPA;+J:3-*#< 
@UQC>.,SS9GZP]O8C/5LB#HI^JQV29MRIH<Y1,;T3/YL 
@+X8=3J$080_ DSTL.N?+49V@>(_EHAL",<JZE=;_G04 
@"M 7'2>\:M(JOM,&8>A+1-0Q[4*(B5T>L84U?3?.JU4 
@Y>(0K\+ 9I58QU.*D8,J_M!0F;4F!%72-W?(#"*%;8( 
@KXOXWFWFB^IK-&*F("JGGMP@T#L3OV@%TEM+5=7>/ZL 
@N!I2C-JXWH;-^W3+U9QQIA!<Y,@A."N -$M:Z72&]D, 
@'9+\U,SU[5]=M2UW-36BA%?:Y=%@T @SEO,3GVOBW@  
@[0*&*T&ZXX=$"U+M.PHETH6FB22?;=VMA 4TB#I;)!H 
@6@.W.,)07+M&.'-LO4.GQ":P"G7N H8L5EK7*/'F.*4 
@J.L+*S+(43M$]+T]AV^U'!D! SN=E&=93@*]0BW5N;H 
@SSC)NYAY.#E (,HYLN%H-'E@Z;W2&?GK!S_A:Z3S*DX 
@/Y,$2<%PGLHI:D+(0I-)S681W43-<, 89AS$6[D%_[4 
@1J%!^5$9K90(8?BA'2P-Z4<*24_NX7#HX<S>0+YE:=0 
@K'8ZY,JM*^Z9RYY6)?,)$]&[H'^ [<3=,)(TOQY+-R4 
@R+9%+_FPTV=:)H =J=#I[XD,\<VQ_?Q):C1/%=AO5-T 
@:NLWF*>+T36Z-]2?LR&AU'(<'A&B*]9QUZR'+]'"9 , 
@U--XTY.E2!5SONGX5S#\6]K08VYV=5&)])XJOO-899  
@+B+(YRN^C[7;-P=NQB&@2-@M13O,IQ J[?_V]!860?8 
@*6E../NY##?FJ+1=S^CDZ[S(OYG^N D>G<$4G%1M,F( 
@$)+6"&[<Q G^K@?,7DWNW>RG4?I@TSYF#Z;^;S:C /\ 
@,(4M@A,6K@*Z$.X'0"K*K/<P9=MH%9#\+J[KBLPY?L  
@([C./V0+CTQ?IA$<8><][H'*5.DK+/!C<J^*2)B8\N  
@P#D:#)M,L+X3C$$ZE@B$$)(J;VUEJNSZ04KPN"J:ANH 
@0.C]^+$>7</ *Y2\T*H#;&B1W!:+?L<%A, )$B!9A2$ 
@/H OE-K:IDPKDQ;^L&J+SFD+&UTB0Q@8E)2F;E@CV:T 
@%EA:_6C.=819/7LJ'[J<%2%1F#_R<D@;F0N92>7B(]X 
@ IB@S8"Q#;=>"26\"39>-]12O<E<WK24+$H1CQ.M[ T 
@46YG_"I"G:Z+>ZKHQ,I!(##\:5\WP@CK<6H5E/D"SR0 
@*X9"TM!6L')X]5V<*U7,$SZ$T0!88)$FH*_H]XH#:8D 
@UJ#@:^Q0^ZU%GO%175 /?X=F%)K6+SW-I>CJBO5O4&X 
@V3%D3B[J>],7G.LGP:,@9G9UKI))UC:?E&;WC60V00$ 
@I#09?AQ5BX1L$5D#$9ISVP)1V(YLT7D-X-X$(>HY"\\ 
@N,W85"NSK'+$[86Z)NKL^3=5&$*R15C2P[W>#A6Z>/< 
@M4"L(;RW]/"DOQK3T5@5!A)S",0VB07G'G K8.\H7B8 
@;6'O.6WT[J8EIXGW+=[FDS'$!F<@D9*$.5:!X]^3BA$ 
@N-;38 E.J0E.-9N!W_%T3$L/\I8;UFK'239ZOVKMQ#4 
@W2S/2,A__<*895O,0PX$LHV,5+?-@830KY^X]JC4X!< 
@=2R?G@I]M;RX:UB]-MXHCCM^5S&16U^ N@U\^B4(;$$ 
@T.F&/EG$QXO[O@&?MY!*1=O#/P,I#C*&'/6 I"9FY 4 
@9^_#'Z5P&V?Q+ISM!@)+ZRA3 ?4'-4X/_<1-7M.(31, 
@#<'F-P[NC5(0J>2"_Q>H.5S^QBK9.D/@=^T?F'IL4M, 
@**I")8-K,3^+"#$6B6)UZ#S6 FW:1U.?V^LI9E5E)C8 
@CK6X-S%F9N]A])8UA<4UBS>W\J2-;'L@YD1=$"=CS4< 
@I&C0WY[NU7Q@16' N!,E3ET5NDI1XJN@Z&LIFP-K.3L 
@PUD4 RAL8 !B D<(2!SYCN#TD504NYHB^KSZ/G.:].( 
@+7KY@=8[3QWTH$N@I8!%C;K]*Z,+^:6KVOP3\Y](#A  
@ H&%>F3&)RUJ<Q0"UD(V"X?#04&Q#0@ITXL+22W.7PX 
@P2*?,L1B%T5K5[!TJQ'PMRLKQ.XC'":S9L)3J)9MF3P 
@82197T^2^SP;W'U 67DV.5-$38(+ 3$;>E]Q$P$?LHL 
@%DXCTWY7CWH,A/#HC7T](0QSPYQ#M*2B-?*<.*6SFO  
@?(0%?IQOA%L/)[\&$R?Q\TC79+[9"%Q<$AL A3G?8HX 
@SG1M3G-$1^N;?\-O,:]#5HAW2$0YK@*W-'K^R,CZMI4 
@)L;'6)K3V[/_5E2TE)MD?Z$@M6:G!$<7<"OTB>Y%/<  
@@R-1(E3-SM(0G,1&P)0XUB26QA_?0A/9JQ7&I5=L_$D 
@L- (\-MWH2)L5_A])2*?4$#'I/L""E/51*(6[J/152D 
@RO;LY:%:>*(;5218F:KGS=:PTU<NI$\AT9TXB,#62OX 
@]RLK<W49HE*2ZJ4%#3E1J<7A39(H:WS!YN9V9:<>(DT 
@L 'Z^0_R5T1UR8<<@HZ)#NC0;1^[E,E"QQ[6*57L!FP 
@OR]/REX1W4ZH17Y]L,*!E&GA1=@O&R-K['XE2.Z*[1@ 
@PE3MILCIK@(J3Y?N;T;ZOA\Y5QHM"VZXH&#SH258?1L 
@C62 /KQZ]<"T;T4#5 7G;IHFIZZ%I*9)]<OO[Y&1PN@ 
@.14_;,Q59(RG-4+.G,>0;'-D(;W17CL37>^$'A*C;%\ 
@[&,V,FEI-RUO*)\S1*3L=;? ;5%9?#_:'/[#J4>M)@( 
@U4SH*Y)5N@Q*8_1.D&O@5 "@3^+]M =E#]TA$=E:EC\ 
@<.F,H"-?T%8JLLX.9I2__,I59FW?L.O3)"ZX2+S">H< 
@^;@6[CXBW$,54/W=XH*<34F[.:?UP@D,32]&X*=7QE< 
@Q]:C"%?!I7,I(7W7=$^,8N>V>Q/[P,H=N _)Y:V<YRX 
@RFNMN)H4M>(2GF2KCD#+7$4? O%>)K=F1VH/9)BJI"X 
@TYW/:09&(!<^D^2-,-&"X]/2#GZFTE_1ZQP&-<\8(JT 
@$,ZS80Z(QT-(4V1#/[_W%54#UPYNZOL<GML'X!T;@J$ 
@P?^80<)6NN> &P!WG@A*,X^.KVTK(1:)QP%VC1A5/*@ 
@TNS&G_SZFW23 $P"=JO3?_0(WB>E:CKH&9=_9+!HB-( 
@JEL>:_XK-&.%5XG%/63U=>AS+R":;MRJPX]FQG"#!+  
@#BV).U#XB"NS%G;2>!MHG-?IN%\+BQ=T:3GY]FHQ(S0 
@KB/V/>U [#_/H^H.%H8 OE'#XKZ)?9K[J_W#>ES7 5< 
@B06%KKM4/R W[QWB,E>PB:U.@TYXBD8&^CQ:(!">1HD 
@$A8:@*8$!<2>7>6+I,BC8WZ44%]X]]RGE"C5NVW4U-L 
@(5T>\U6ZP"H-P(/&#\9?KT_X&/?K1V^"WF,!N.;.O<4 
@#GXJB-=GU\Y -])]SJA?VE5O/P_33?&S0&K2<& S02\ 
@<IFT+ M0DM3^1O. IY\")J]#P@V?"NC(1WEA&(97[ $ 
@S&EGU,<X*K()8Z5U/'^:E.B=258V)R'4XT5&0CECS)$ 
@@=RXHS;*#2'WME3VN64+C-S<\"@ P\=FY%+"(=9?YTT 
@:$H<%S_ TQ2LS U(N(:-FSDWR(<K<%S:A9;QID>=(:\ 
@E')LH4(GS/F%.T,Z7^&D5,E>MPEP!$@]*1O<) 4X-;  
@,O1+/#H0</R%9A-EM[+C8BF@^HS^I+)@QB9K"DU)ZHX 
@A9%Z8>\A0*M_BAZ?N[V%+.#D&UI,>N.LBZN!\E=GLOD 
@4LHOQ:C)KVL!/O_I(9@C/@CEU8).H3K"0K)1(,\0O)P 
@X<IM2#G1>\R1J\G#,L[YMSADR$NRKE>M^)_!K!LXT58 
@AE<];Y;@=4<!&FR1R.1$6$D#C__W.+4+:RG7]3?J[RH 
@]Q)58[0N=+D>^):79EP'W'4?,B4E(+X'HFQ#ZZPZQY$ 
@Q5Z;VU#!GTMC ,?LBQE9";CU:BX<Q6(^VL?33T9NP/< 
@2TX^GQD*3(:'8#55E6Q\G/+FAR4*J.%K23DFH6D*3BL 
@'(]YV%)O7%CY>N\RZ]S'R=3/EV'&7#NAP-4C">(Y".P 
@,/&A%+MH8]*@5S0!5GH#/6:U0QL1\E9TX)+JR99@E), 
@8=7SZ& \D4S$?N5D'Z<01()4\EP4)\?[=*8,3VL?J/H 
@BX10XWPFW86A:8^2MPDLY7/]2 =GF#S6TYRJ=$:E$A$ 
@7;)S4+<XZ=7S6,CQK8ILZ?D%3@W\H+;H%MV'[6-H![P 
@Z?93Y!W/ "1_]O(B)/ZY^$4RS,=*1GM3,[@VK#H?H$T 
@6\CDLJE7>"+$:N$#>[ZU12(*4JCZ=B)P9.HY_*+%EU, 
@L%VB,NB7*;.7(M^@/462$:\?Q4/'NC.N5FZ:BTN[R4$ 
@%A3Z7?7/!:!0N"S).6<Y2(([IM?;HH'P\6?>UHBJ+R$ 
@&:%J?M<QJU5:(WC@\D>8II0R%#&!A@[NIFG__WGM3U< 
@6_ZA3X%&.^LDALUD[2Z2>/RWLM0W)38Z9J:M$IW9'X  
@%R]\W:G?EUKV-\4_<"-RLQ=@Z.<('A=S-WE1K]G9D'P 
@F*_X^]/:%1W*_@A*0>B4HF"D\7\U/RD>R8C;MOA#ZZL 
@7R.%<.5>=? G!;491,2>'4*P[.*MYQ+)HOY^$P>LK)$ 
@#H>VRKUEP4'(']X(6;YO %ZD Z+-B^/VFLM]\**("S$ 
@:VI]E9Q::TZ1,LLE.,O"S+G=,I)82PL_%N"LG#VTL"D 
@?)H2.:[W!(K)U_-]A1W'6\(FQI XY)N(T*L%D:?J1'L 
@Q!80&J/2YT(%0E\^^AIM&'@I1!AE>[D)@7&'B;2WVLL 
@L^\J0W1$8/ZX#/N'M#Y]5ZE1S,/B[&_TJ(2-=)M]$$L 
@=:VAMTN;\XPT9QV@#,70O%,2YD+?=_[8!_21S+NEV 8 
@I:Q/051K:N65Z!?-Z%N-DUX*6A[AUR3;$=H+>A)Z_R4 
@,/ %2KO0+;$'OII\SP1O_.VB6ZSOD,R3.N43$99G1!, 
@UT3]HB>@/;N;*4.ZTZ_5@\=V+,M;]7F(_*]VN*Z5C!D 
@)/Y<)D*LT2?:G''6X*B9W"...1Z*D1[IGE"+##JR,-H 
@:_,9WV%=X/&?1A8\C L\YVJ!MF$3!;(AMV^P\+Y[:6X 
@Q764*XMLY85H4>]AKP7K.E-;7@(C&@FPQV_DW6WU4F@ 
@D/V'@,Z=XG^Z:9F]8!&P,,'6/G"2V!..SVOS_ ?)X$@ 
@^JYC4)O!U3C <N3)0'UYUQO(^7GA=,FG98$3FH_%7)@ 
@UVU6[X& %TE-"DC=G?P<=K45"+[@;B70O]-%RA+*F(8 
@0^$E8>KCUL_C(,QF)]A^3;E:D0[@-:"MMDW]60G*F.$ 
@G?A80P-,]1269#.1/&B^01Q/%7-#1!NW?:H^V+(BAGT 
@."F *Q.O/)-AMJH/9FZ;-<F!55N&)*L)[ E'[R/?F^X 
@1I\7?8F&TE]R"^HM9HD#X!;XD;'2558MV9EMNC JL!8 
@86?SD.SK%BR#3B=U^(;:#:J\J#$EM"L0@-CET@QQE'0 
@YA\L"#:"B\FC:3C8@-Q',:H%I>HTDU"8? HH]8.O Z\ 
@GWS!LJN?EK UZH['$B](>,NY-Q#AA-.C<0(;2I[E+^H 
@6QKBG[ IF+*\KE<)#SVIL&9T$*4G@Q6>E%+F,22*O9L 
@_=;+OU%28M")[=,M"6^X90VZHAY,4*-C?#2EJNWON^$ 
@]$BIC]7"]2$K:A?*?;!SG#TI;).SYIN879RL]A(8)!L 
@AA ,4@!P1DLJQ_OO*$YB#>UY%:;JOX$PL61Y&T'<]L< 
@E+'&#B"N?6)ZU6[SDL8H<5;I]&<2=9-%)0"T)F$F[A( 
@?[4GBDX.6G4>@J\'_BB5TA.B#,3'DQ0^*C&.M5R#N"  
@4+EM93\$;Z*+C-O!VM\NG*( C'-!+-0<]B;B.YE*+CH 
@*T\)]#)^3QK<#9FN+,9^PUVY_Y(J6Q&<]VQ,G/]=YMT 
@0R^BCC8*$ODA4)[X)9B\%2&\G5W3-G!ZS+)-DC+2Q;, 
@<KJ[07BX18K8I(2\ &&F37;W^R2%+'"[B+#Y7J3DRM8 
@\ PH*;3"7YM)C0&O^(<E.F<4AFE(;UN49&P*E.50U@( 
@> *4+JD"]<N\F/!A53HY8/L$1_X5*-TI9$,4V]X8BJL 
@"O5=O%UOA$+@ \P$;"P*K&)KVPL>Z?*;:[_X.!Q'S.  
@%",]*&^F?2-'3Z/=*P^(#ZS9KS5_^?%9DMQ 6_=IG < 
@[),=R KCO7@25J0]]LOQH@$J')%95"QK1R*]:*I(24  
@LDCA*TY2FN9,L+>S+[4"+%-6^AI?/*L:9G&J[M4GR(H 
@XZ\U='1.IVY5[\>[&,\D7[$6S2>TOI.'90R[ ] <71, 
@R)99FHG<SMP0#"O3/OSE+-@K@*]P@Y&=XI) -PP]0+( 
@7Y>-CV(2T43+7,.6'QL:8,F+6__K0:YU"=B&_?Y -T( 
@=(Z8.?D/3Q_XU21 !\X XHJS89.!1UR1P_&H=NZM/-< 
@Y[$[7WDC2MU=GL;&Z[IN[8Y8!\,O/PEN'\(,ETPP!<H 
@SZN5:PGV]0Z*&3JIV,< 0IHIY%U93TT_E/+B0#W<W.T 
@ZJ-\P/#-"L9@AL=K;55MGI*4!N#VOW3BI<HF5?<] "4 
@?M;6",GR[.IKYIOQ"[@(W1ML8JTVC]CSPLDGQF[D!WL 
@Y/Y!#6]63$7I;JO;2YE-PE*BH_PUY!C^5KC;)ZAE+:0 
@>5[-)]@!]TY.P@+X]/](#4+#\;#:.">&CTEW =;,#/\ 
@?8B4KK),%"B=8@&F+T#UFQ3OU$ET;[!X2QEW 7\M+^T 
@NU<*:B3^G$,.?%Y#*R^DRCX2QJ2ECKSP ^*VI=I2:2T 
@98)6.6D-O=JBI2R<7*UK\.,,K),RR;=V99>=C \B^KP 
@VS'>O =.ADXH'@BVW*N$Q*"M($XTU2M*]B;J"E,V=KT 
@ML<B;IQ_Z*]@&!(\SRQBHX]^.^+%VQ3T&GYM^:"Z2QX 
@"^C5RO"HJ2G.-ECR]XT]XJ"[:S@<N JFL";,FI"W%W, 
@\EA67ZC5PE@+E5KQB2D_OB-8?#GDC1-H0ZY.PD:']_$ 
@1M/_KM*+7)=71PJA@I,/XD"PA$XW.15V?=]X$#&A1P4 
@F5)$4,+(S#'3E<RQT?F",>D"L05#+K6IY2BB/Y5&5'  
@P]&]#NPD5WSO?F]@DB_Z#>A-2+VZO<D1&]0E$Z)Y5/0 
@\K<:;(*CGHC]4]X$/,8E-<)Z\KJ/6_$+9HC >+)%!@\ 
@V&T#8+<<;%]FDOBTW6KF$Q XT/-+?(P]BL0ID9^B@W4 
@7^B*C+]K0T_+X:!%3Q(SFF3.0$S/6(JQ7$=Y!\:^,M( 
@TRUM4&#AK@I_FIFXEPQUBFZ3NKVH6J(G#6BN#4O?9&( 
@)ZK]J<G=8U. ',Z(P#A8T<&&6K/^1M-($K_;WHVC1+L 
@_/6KSG"1A7R@*IEF8M78KT< Y0)P3(5$__"WP7-E%/0 
@6HJTS/ 'BF#6\C4*\" =!@5RZ4!=]ABCT!+F<Q0M 3T 
@H80'&0\202;,ZXZ3A4.!7^N1:(HN+?A%#&M%(9FR+TP 
@JT&#RV8)(+H8:S(M6R;X<'+4>GY-?/#NX G<JZP(E2@ 
@O'6#1.UY;;V=-ZR6+ZLCQ,X%G5LX@P^]#<7_SY#Z]D@ 
@7(>7NE*EE.X%]^[:RY++A7T+\'L63J 3J?6.H;HF7Y8 
@G&-E#6(Z@B[U'99?OC22&TLXFWN:DJQICI@7!Z24_Q0 
@@B'([I6T,VRJ?P)CIW-.&W(W;]F"AZ=F78\:72&Y12L 
@/!?5\!0&2-(SA[;0VNE?!M73*OK(WC)>"XH^^"@_HS4 
@4O1"C%S5_9""/<V,E2I>I"UX>%Y#AN*C[^MP^(VNK*L 
@''^J8*8T2[Y?+E4JK'(^]7".=!E:*:;3;2JY?YY; 7, 
@=!G!L.[,[VE7G4NG,M8'&'TC".AFM5=+%V<;9+BL;\T 
@$!@BX)4A?2&;VVS?:/0TEYRNI?;SN-SRRU>T:;($PGL 
@D Q?_/QAA;^<XT35>1$&VGZ#]6*,T9GMZR#SNTTM% L 
@,N!2IZ7K+M-C/U#YF%S)U(=U]4''ALL2W#,:);NP08L 
@Z)Q_WAK(G,U<&5:VCG'?KJ>7":>PU<U8U&2I"^;K/+@ 
@K:L"3)>W>-B=Q.;!.G#R-ETXTCJQE$W!./ND^'X*?(( 
@8HQUMTH+@MLVK;XYHVX:+WSKX:=&@;/VW4-=N4X+78( 
@:MAAU&+-T2&+:&FQR[D2?A]1=.</5W>IO]/'Y.;]KX0 
@2V"(EW0V=+0)_B2RUNT/H=\<9,HY%)!E:WIRAU@R<)\ 
@PA;_^=E!NN@SUE6B4ZA+4?)*]AXY@,Q!IR=#6OW0$DT 
@:U/>7?@J.CIU3EW? Y4<.#_F%TV"LA">051,!K1B[+4 
@3AV.5! 5U3AO"-[4#W.^0+7>:2N67%0NY$%1*SJ.0-@ 
@&N#:T[>T+@U:_.B5=O&^^-R5@O1&.04.3_A_TJ(DK$( 
@<H?)6(XB":MR$9_P+;E<3GAN*-FUJDNDTLJZO5?#_=  
@F7::SJZ^C\Q\'GXX5:L#' VXH>L<H R$4+@V"$]H4FX 
@N''C>R0!)N%OF/V[=;D68>DD6 C[3X^_&=&+R%01)?  
@!H*9C)-EC8G)6NY2P)_IP>E!5ZFM$;0?9-PW23'"ID\ 
@5MC)HWJOW\&Q7#8J$%_(BD6X&<8+^T</WR]<3UHR2Z$ 
@P^X-53G@X\KBPYL$E1B"MM]G?82,ZN\A9+,2HMX<J4T 
@()NT9/0_KSN<TZMM.Q.H_0-@J'7@'C]74%JS:_F?2VT 
@"NX4U@8+V<X2\>[+(&VE)QELJ$.K D=<4,Q*^^6PAW$ 
@YU)-)BG:"+JWGM3W1IY.R 0RW%E(V8'TABK1M?D9 %X 
@&8D$QA@DLIZ_8TAZ;=C\VA,G#-&WIE:EYYS(X9^O,%  
@<PZK+:&NW3CZAQF4Z>FL%<+]TFDB'_(G *]R$V1TKIX 
@LB?@*"Y.8-<):UWMXRVMJ\D?LS0OWTNMXM=LA0Q<G!< 
@Q'I33D9338?3 X.G"--SE?$<?I7U_)SU,VZ#1\E94^0 
@=$]HQ2>"Z 8O[-KF4HJ4> O5&W+XCF&U*T&"2M<PQ"( 
@QR'087H1EH>_#K>9UW(WTMA$>4I*FZD!WJC=1F_36^H 
@-;_Z?ZD]''\3^ME8YV4A/E*TG!07;K=AD\1>?O'^'AD 
@C+B%1K[YG.,NLVLUG?C.ATQIR#(!U"@UB2UZCI0C/X\ 
@!K0J@&_/5&=;^;,70'.0B@[. !)-&+5\)F":P4;<!FH 
@LQ7@>!<X!1J5&J"@023Z%N[,P=*UT,(>H#:.JM,9];P 
@6@4A)V3;2D8/8UG\\>3+P9C"76>R.T\-F1MBAR=O.I$ 
@%BKHH'4KC3*9HA>$8"-.]_!QTX$7: VU:MB93L>K(9$ 
@<;1.W00;G:9_0N.WW"D6!.N_4>$*!%!>=L="]0J_0I0 
@P!>.J^^F"Z+?-IT#0$*E,:UA2F"_,<\C!DW/)M>NJH( 
@J8[AZ%U]C=N8]Z\P%=KE 92(=&=!5."CY2E1PD$"'.H 
@$&8U8(_TT9BSW_%D* S^ROY,(1)(<_TV=%M[792A1H  
@YIFJ8N0&[_2O3ADF+BR79$ ]&F04KBRJ/ [PD8K<0+H 
@N@G4_,B.3,R@T)#41 >P1I.%,IGUCD65IY!AOE6+8XT 
@/;LHJ&T;>\&NZ^V_J7_W#;4+G+61P_,R3(0F <0N\WH 
@@E?TIB+1 (#L$7Q'_F\?(7Y#+\N:WN4Y";;M"-]"D$4 
@GE.<*_4SJ!_=>+I#S\7 0[6D=M;GF\I$@"5X]MD(NL< 
@,T:/(8[]P*J=]=L[ZC)\?447-2R]6M7DK(9#EO<S(#P 
@7\&$8IVS:$8$0;:(YS767#E+W$OXMHO$;T\5O]?Q&3P 
@D*1\WR#JQ)0B8_9[E8^WW+3?(P8_*LQ63,X@5/WJ)YH 
@BS+D:5;P%*UKC<Q^HV\@?5%%U%78NL F1BOC"THU_04 
@ARFH:-DP]N94=UN$2UU@7[D9WTQU8-S:,]R"DT17ID\ 
@L_"0KAF2WFH.ZU2AA4^E<[<D0I +[L<:LH7$%+-I64\ 
@5C^QU.H.$59Y_1/T0O;E;P5__Y9\.6.<F"JIFO$X71P 
@M]8[W^?="Z)'\3GU^6,,V6\Z2K*Q>:<BEYUI.C+AP4T 
@Z^DS\RO$E)FWU&/FY%3,A)?I&&29\RD=ISS>F4$X9@\ 
@%!%3\:%FW*/-]= GQ 1+KWZ^9;5Y=*CSR55$71?LYE@ 
@:O-8,@'T\8L"K<3$ES+(T]5WZF@4M)*G%('&V["WW.X 
@^P9_NI@21A3G(O[H'!RY,^H*OFUQY#V3O]F)'\KK"$$ 
@C\9\M?YS,#$&?G2R[",_!3.2(?7*7.KR,6=BE>VJY"T 
@0AT1@*Q,'E<QF%ZU 'N.]E]:IF5A/!.2PN[T]BK"X \ 
@\-AL@4**G1#8N(L>"2[4O%=)&T+ AMF'6/XLD;AF' X 
@-)]G>MVBS$#X0/.EI&?2(R]:'5$5\]RO@+M?M6GWP/  
@NI2K#=.:L\_$91J@49_^@8/:/O"W3@^VQ4$?;/_@$_H 
@\UHFBV^8]? <6(:"\_4[5(]6-XVR%W?&CY$A3"^!'@$ 
@XXXWVFUBLV)]^I."T671\BNG/V(GMV^"P"HH\H@N89D 
@WV+@Z=";"&J;J->M&U90K:F"_I14A >EC&4'8$]#K!$ 
@RK97B%G$J$[XXJTVKF=(D]B6M9YV<M>B4&U6>G6B-B$ 
@1$]DN3I@/I+4E^_"5K&PY.FJ^RO6K&:TO ]V70_M<4$ 
@*]C058\?B:W9JMYW-O502I@^":H"&"NY)ZEK#$53I20 
@=T2*SX.A5K2[TYQXZ2)G8:R378_Z94R#01L\9"+2J&T 
@>9;&&#F@KA?W%2(_RWN!=XTU5;U+7H9Z.Q<#,X>YKX  
@]9Q2,$[\#FA"O"[-E.(+8+SQOA*HIXGW'70O,,#;$%, 
@]0N;^4$F]8[,4?=\>Y"D.>2R4-4F2W!#886.IRG?SO  
@:B0%=.W8#XFR12P@\H9NA3>!M,)SJH1A=]N#";^+WP( 
@#"C %2]GV<RL(@9>AM]/)&H3. =.<666!!T=3(B&W<P 
@@AHN>0_IX5@=>PIZB%;T]?Q-R)"UZU<7<?9<ZR>I]/\ 
@F(,IT'&4H'A3X'</H0NNY[1]^M%_1TSYA!OY8B6R'N< 
@A)S0++DHP+75-:'/<S&0_]93<UBQ(E;B"HQ9$*?%I,P 
@+@HVQ@<6J+,*T(5'B:<M1V<^6*UMT<<!B)!SX33XQ/, 
@EB)DMO /)/V:[W)#[BD8>AS5<,HW*_D&.K(?E7)F2MP 
@H7[\+B2+01:+.4?8!D(/'?EI&NOL21]5E:G_5+\*Z/X 
@3YV>>2G;!*\%TKZ;97V0YDE6#<^R.")5DPVS"OY.-8L 
@OVF9,W051VF*#&0T\Z:@%T98\"25:9@>7N9"DP"A4#P 
@7608)^#Z=_>!M,&L##M,IFH>,A1B]W>+.05\UP)[ZWT 
@A=T++":L>L>YK;CC.Y.4YQ88=F+?A^7.:P[$0#3-I5H 
@,\>KS%GJ.G:(:<PS=-O445$!0VOLP?D5XW[$4!AP84P 
@4BMSC;?1.V5@+03IS-$FQ<8&9L)?"TM.74:ET$+T5[\ 
@4%TQ>F_T$OK_."C8TE/&VZO66G7J5E"0(4E.'_W/K:D 
@&M0ZZ=\K%<,[Q>51E"Z,1[VF,PFYQ,V6G33?$R?>A%@ 
@L6<'8]X(+8$V.<8CK')%EQ=B]J(8 5CO@MXY1$):V'P 
@7<G"* CLP/V#JL:17)[Q,$N?DFSURA(AKB7+M_[4$;< 
@H"T3D @#Z+,JH0@[&S]F(".Z?)GHU7 $+C1#V?(55,< 
@E<GA&?-N/]N_96I+.P /X^P<V,2 +0$'WMF5FO8<Q54 
@T:)H-BG$6M& @755Q&;1/78Q9&&-,&;.3%++1P=!"+X 
@->G?T[$C(B1?*AQPO?643SJ]&&FF%GVU:#Z,A;35:S  
@R[[45^8VV:8Z$8- 3I G",=8_??=.31/J/.QA[4M#<@ 
@0MC7VO;N/[(?A;RN";U#?-VS/OCNAK G$=+\QTV^;DP 
@4-^KGU=1M"L;MU< "J%>WZ:_H1\H@7;SOT?N895@X6L 
@G'0DQUO5_\*5.C++!'E-*RR>PD4<T$K[F%TM\<HAZT4 
@,4(]C)#IO*6$6B*'HY)?ET'K(/3/JXE0/:!Y2 H?;*$ 
@V%]290;"$ZM<XC'QY@_:16[=_A]CY4T#*AK<5\LQ<NP 
@T>/*"T=A:1KO!D<U:^.?CT4H$_HG5S*[X(%+WK<CKY@ 
@MC\/5>C14, X[@=)\2'%K@#1.]F7F#%MCK/U]HM-XA0 
@M?GM'F<,-R!ZQLJ4%,,"V1#)%N84V2D!(WO%],XK# 8 
@!X$#=:AV>IZ$$D[Y%8#FO+-P?\B+$OU19^,JH;' -?( 
@,;*1B_,G>7X6="%3UJ-&G-<5I;1!B0J&D(\#EIZ(5%@ 
@T%%=Y,$6M?"%<=GM"6RP*N!\-DOWF(S+NJ#".(!-S_0 
@4SJRU<ZG=],%L6/Y-24!I:?DIK?BS=(X:-J=MW1\I)L 
@9/M&?M8ZZI:1!("O08"8'KN6C!T^LUV"T>6++B?^:E( 
@G@HE$Y6_LU T>Y'0OZ/T-"\#IR@47!&Y GN^2>PY5%@ 
@.%_+WW FJL::PGT)S]D-6*_P;+:O?'W(F8H&09.*3?H 
@/"V%7T>*L.!.AUN^9AEC=VBP9^]IAJ)'UYI#P72AMI< 
@=37(]6'-K5#BZ8D@KO09=35@D9 6;_HP6UP^QE,2<DL 
@Y7QAKJ:JI]WOD_]R@3GCF9XWMZ>QZV49QFT'/HFC\.  
@6 3A^CHGE_!3>(^N.J$EH[_#%:VC8[("#74SO?"D:D( 
@S74T=O3$F2X+(5%-8_#T(MMT7D=I[NF;FY8DET;\G/$ 
@F]E(:IGS*&OO2BG._8F&))IVLP-P[<D2WV9!=CO>1)0 
@C,94=9N!)[^=KU$\1 _ET"]BMXNXOMIS&0WRVQ62"$D 
@Q$S#0"JG$-#/-9D^B3ZTN2Z8?0_HP9*-DI%0?]"XSE0 
@M!B O8N^N*;R$W1O]R)GG![HB4$=Y94$DXWP,S:Z<L( 
@W5-2#O]2B[<K=TEE$9F9"VOW )1/IY_$G.L9")!J](D 
@3&O21#QID5"LOC3L,C:T!NZD8GG:-E2VT^Y+?)[=+9\ 
@]3TIX,M_\"Q#3LE#+O@[NQW>E*1R@^H*>H]*J& #MV< 
@'DU]@'1;.EQTP5BYQ?VWE,"\P+QVE,EG?@8>JD#FP$$ 
@W?V2UD?S!_^? W:H/'?&7](E.RH '9/981"H!B@$>5( 
@MI;+4"PYW5B)[00V5%LRKC_FA/2?PL#!86JT"DEW^,T 
@GT7')/\(LA"3SD5#I\4&2>/B=6A=8&2J)M]QVTT+0%< 
@P/&ZJ5-D37^@:=&NNOI/8:<H5EN"1V=MNSFR?.@0T(8 
@$(0":J5V]!#!PP'CSC.<WR]&D /'&W8^TQ/5(CS$66@ 
@5II,D8FF03UA4YZ!T-_TG2.'7V:)!Q'U(:XS&6/F>/< 
@O!;>/2@@+LX@F/XA0'F*&_YU3W:EM$6=1I:#E=Y, A  
@-8"3W9BB3]E>7'#JNV._MG: I4848>!6^,"@ B0V"Z\ 
@F0[;.@^>=3,#K=+A[2FI4$CFV74JW[>2^$/09M#B)_P 
@/<P!J_G8D(H=X&@JL2?E.2)2XL<JCM8 WX\86:);QW@ 
@9P 1$Z;W7W[1'TDB[#X%R\8317N2=IT[<.((UE),R,T 
@!K4CBC5M6ODG57IP-@?XIS'\=Y]4^*&HQ&.FV)RHEAH 
@'O&(?"]OWMN,'"(CSO:W7!QLI=\@QY2.-'$_>+("P(  
@JY,CZ@E-CFD<"H/F&=!T;&7[7R]HM6>[Y S@C 6ZF$@ 
@H@RB-WB%#^LJ$XV$C#Y,6%_:;RL_H8J_#L$GM%3Q !, 
@@XJK W[5'CG0]L6U97I86:%S#7\['%%S#>397;NJT[P 
@GUB]L8R$)D'VMFVR:B!8%:U;2Y'6C:HAWB[3>\V&#\$ 
@ZNPENH%E+_G<CV=7N+A>RQR;J7Q6?:.0U0&6Q= WI1@ 
@\(U>K6 ,UGW*+KEBTA#&)_O[^R5UINL*^8CMDH%R%_H 
@^G_85RR>?);V07I"A:O,NV)@<XP[!TU%1OS>0$D4.%< 
@Y>*0_T"<&,(SB\K/@?%87T&W&NM7X&;3??&XY@2_7)\ 
@F'\8LXFCH/BI$NM;20JSIOM]\T8-@%,<TB/?\^?!#MH 
@*A*90,_HB.C%)@>36&VB6VM"2SE_A63+=0P.2ZBV!U  
@CLB"HHIE4<%M311QX&!K]@+-DP"=[&#D!]7<8"2=B*$ 
@(&KBC7OJ/4#Z )8QF"$Z#L.?I+DWL$S>=N\9WADV_NT 
@H G\UE?%#&0_(!G_CCU1(5^$!B)8"4-I^7P2@Y4N_Q\ 
@Y]88"QSS$9SRC&^"3#F6<Z7,&G46!*$&&#^^^H\'K<  
@A)(1L!C$#[#))C#Q-*DV'7?V\E\Y@C\$DT/!F0Q\ZXT 
@AW(W-Z^T GEA"+MR9CUOC8PJ&H*;XVE[>C:^4,!K$B@ 
@)CGAM=4<#A%V]%+3T83N-ZD,/G+.(1HNI)&D6.1BB\8 
@53YZM:2FK1PE:ZNQD5N4XV:W41EGG22[RIC7)8P'\!$ 
@K/^P>><&WL$^;=)\\-^ 3#V!OQT1JD[3D&K3H-BH &0 
@%V<&(1>=+?#OJ?C9YP64^K]ER>(E,5(<>C+$W*T()BX 
@(9=6+6GX5B5(\R'2I_:T<\=Z'&E$"4QV<2.#Z"II&-T 
@5!#4?H*B8Z/B<!GP!-XMJK0T+ $.N-I4X5I^534]Z;( 
@B/W%T;&>*@8YE]TRTUEZH1^OCW@/&R,^0+3'@A-PB'L 
@2<5NDH,2JII(5X&.(&OIR"HP=Y#D)?8F_%H5W)TX6KT 
@[]<ASBQ1WB)]) K"<?F*X73&"@0)G6[1@6*XQYT"2N0 
@S8D&S8'^G/+ )>JPG0>)QVS2L& 5)?[' G;J/W@LNR( 
@#"TJ7_O*DSIU:HKO:N@F-KP\75TQ[P@=SUQ0I+L9W*$ 
@A/E<F[*W-12O;HBSC)^Q9DFD7:C) \WN<XTON [DR(L 
@5D(=@-H9#^4*?,[A,2J%_H;^DA&QNH<[?T7_B@*_A#H 
@2GDO"] 0\O1YQW!G2T2S?A+(T:O0&:KK$CE 'A%B]4X 
@!Z60)9YM5*J+&_S)"E[16&F$$;E N:E?O&<IWU693_P 
@"/_5OGSG^W<QX>\800D_N']G!%*QRMSLFVJ4#I(HHY\ 
@__8,J/0B]I2E:Q(C/T-]*O;F%#23'IB0+RC9 B(\>-H 
@<VER4W5YY%Y]V(1*=SP3'-2-Q4UN#!2Z+-!^93#O0)  
@QV.T7/Z@R3ULMTJS[ZNNOWMZ44K2TEUG.Y=3+3\@F50 
@DTI:*X6M^ 92F94!'P/L)(N[1/=:,SX-?"RUZ#"AI7L 
@VZ@VU?6Q 2!G![_L-+N@$X9NZ  ;T3<52<O\@2\^\50 
@E<Y3QO<! $2*Z"X'1B%GWC:U+@J^WL0&%OZF6.@K4L$ 
@B'DA4IK^O,VZK5V,^/(,4]->Z*VR;@RN$YJD30%?#%, 
@V-Q>$2H&&)#KHBP\#)F6_R.W&$&7YM#2M/:ZQR[S">, 
@31%:I@0)5Z^!;!69D40VTO^+#(]!CU#*#]OVSNY#+ 4 
@FZV=WQVT")B^\E*:\6I\TW3H+>2YPI3*X&%I(-Z26[X 
@ZY$@P$\82>P?: TDSDIW+WK.R4"<+IT6[W<VE@Q_+Y8 
@)-6*8NEIB@;QNM>EUA]\;Z$F;ORSJXGPL/+#%1=[C\0 
@7&YSDHMT=^:JT?K#P^EJ7>H-&=PK)<-(TII4B64\R7$ 
@]R>*Y#@+#404<!R]*P^>9,/:D-A<'V*%G,22L8!Q&A8 
@#6ZL#:H/PTUB(X6NF788(F$18=U#N5"/H3B&Y%*D0\8 
@79=F'ZH@>2X!1[#QSREEQ.,J\P\I4T.BVNY"6304!60 
@*^5$1H$?1&MKN#UC->3RC+@A0S6&^P\R"]82>H<<YW( 
@7FL/IE_V33&.N1?Q0[1;Y&S+A.P=VD(::;A%B$ONT;D 
@PW8IW_Q+$VNQ UQ$Y6[NVL&WC:T..&W61!XLD:>?-T4 
@3\BDXO>(!K,^PH<;X;XD'[TQ-D:4?..%,'QQBZ9\2/  
@\"1^/S'+1UU6!MX('V\G>9H)+\\3"!I30=FP' +;X:X 
@QT#R7-%6KG<P24ZF<]$>'M"EFJ\;"ZRUF:^TJ')YQ+4 
@MD\M=5*KQ X.%?<TSG#I=YM0N1GVBHQZ4+$EMN?7GL@ 
@V.)L=5WA6A2P'=02"?$1CD!LO'V]8/ZW]R,FP1K\4YP 
@)A%6PZLJ0@K$6T<\->3<[B[&Q;E/)"U12^8<]=4F?.  
@4TW;YJX>36+->O@G<V2,*,=OBE@D$=PA\-XOI5[%A#  
@!JYI'19].,"45#19,1N,,Y?1J?[NUTQ9-N!=^^KZJ1< 
@PPAH'S WCG0#F%=&99I^]+5$AT&>.G+CLI=#/"G63L  
@/BEL^.:?KF_TW\S4;AED \I"3W.@$K81[F"-.D5]B^4 
@NFDLWU-1)21+KLK*0^)SMYGO?6U&:7W6>VDZ!'Q-!H< 
@#+RZZOK^EK>W$<VVP=<#KN\L5(-_MC92R#<N@0?LAE, 
@[64#6==R&6/3Q<P8^, >WDX'7#%Q[SO5<#;#;4[=_YX 
@6^-G!?.J!6 G"&+6,4'/5\S8I(J23^2I4R2$Q-B>U/4 
@A2(5,KG)8OFL_\-.,*/ ]"5NC8^B(3:=.1M!'N<A M$ 
@C>#A-A <-CQ:![(*)] ^I"8KB_..J%+=Q^UB(@8V#IL 
@_M))Z5I".L/)( OX>\,#28Y#1,YFKX:4$Y#=Y*%V+8\ 
@3+C&.MT!HA_AUYSIU3'&!$R[!>.5^%2-+4=#93\N] , 
@OK$A1D-V!0R'XTW9[E^EX/<R@8*G4!E'3)@2..5F#N8 
@"JE9Y"2FE 6)=^CR3C;-F_<(]N?Y3\W@(JD%SP4[W%H 
@,9E.^+_8_T.RRL.H$.J3<&9F7P'Q&\.*??A^'Y>TK_\ 
@2ZLG< 3" ;&9)OY@IYV7?HX3P?+IV#]MJX0+6Y;I/!T 
@+G@CFF5JMMRII"2$(K_(9F,=2&].$O@EH?7%C^+Z:)L 
@A-XV!"OE"U6!A1GOMRNM0B,.-5+H->I)C9M,O!C^>?\ 
@3/2+@&=C@74I9<"8;.JL=A\V'!&I 0$Q%-]]%^R5"YP 
@=N>Z=*Z3R&9=3&P]LA'70H/Q;?-P>OB0_Z[6QD6\6A@ 
@IN]GI>SPKHV[JD/)I/^M4BNJIC7CP0VE^/[=5L.IX;L 
@W/32X!WT5$L[-YZYEX KVU$6[WO,_TU0I(#]ZI$91$T 
@P%H7<6_G\JB1O'Z6Q@P52#M!/ <1.D9A8 [L8HP,79P 
@__# ,-L;D/>8(?IZ('I'?Y:>T7BK3QY*SBUPI&,98=< 
@@0/#=YB:)1:KILGBQ-L7?[+189VA@U\IA<%.%^/XSV8 
@7/& BI4X0[G.=Y;?V\9?X G^_,$;GA[-Q*AOQI  SW\ 
@ _(*A*B&T.+!H#QF?M@'O[BXW*G:YRV%<#52></C6F\ 
@@^]9M6M-@*LSC4$MS@ZBE@TM]N^%MQ?FQT1H0#-%6M@ 
@K/";9;Y'JC7+?3.][OI&>;$F.MY?$3K@>;^;.Y<=L;X 
@="?'DP@8>;=>AX6S:?4![KLE%2[15U3UXR YS7W.>LL 
@[BU ?_7?G=HP#'P)%"R*B%2Q[%VX,:Z&)JRO8B#4=WH 
@W.LB@L*3Z\AA_CW<0#A-;HR>C)+K2I8PC$\RFDQ/V[H 
@<] ]1M"F1@MXJIG)3LO!WJ^^K+"!R%A4VUGUDP_&WH< 
@!$K*]I:S#GB1/>,.3ZPX#_W$:L21\<?)C;71V-Y"7M, 
@7O\H$7OO]  M&2F@93Q(#?QL)0JK+A2LO1Y(9+(?&*\ 
@J%*74G7%M:*VR9=KPG9%01@/59NW!M..G%QMQM2>$$T 
@.;<1/T/L$><TTE?W@?&!%')2HJWB)FM;E(9V7);TBVH 
@T:79UK'5SFZA$GM/]0*,*UIK_T_Y;)MIK_,"9!A9Z"4 
@.%MJB:0"Y69/=@J>W523RTA>K_0/$JF,;2)II U7\]0 
@C':-6?E_@2.*]_4[H[($Y]M)Q[1&$/F'(KXG;]<-OFT 
@)ALI&+N!W9&7'1_!)EU&[;@DDS"GH@3%KZ?W;@55']< 
@>FM\M) %Q[&#NVN2&ESE4";X#IYB_91G.TN4),,NMG< 
@);+.C15(#4,[[-A="&E,6-*[F$V!<<.\/WRP>1K>'H0 
@OU9%6CBR YS.F8-0#U>6_FOV;4#>!(3LW\+Z6G.?$P< 
@9AD"Q_+BVPC:[TO&J#^]ZI^8KP!_'X8FSB'I$]E3$%H 
@+3? PF.#9=N6LNB8[!#IQ(%[T#:F@@8 S]\\C7'.6%( 
@-@* CN1*DWP,JQN2Q]^VLF$'OK_NO3LB.NJ+A\3QR.( 
@!$[+D$OHT'X& CP/4&#G"G@[P3Y5L1(3DY77B6"J_K, 
@J:K1TGL ]-?G:?3,VN2FU6[L .=>W-K-8N,1 I?BFJ@ 
@Y;__]HT@\L7^/*#U;\&:I=%N/Y:X:#537CT:DTW[-S4 
@?FG9"2>^:/2<KQ'43_318,W'2$C0'/'V;15/,D0%FJ< 
@^T\)68)CG'L"DN+P-<7G,A<0C)/SG#95BM=H5F9%;X4 
@W= X_,6/Q)TWA8\$SI.TV277,>B:N ,L-SXFYO]!@&H 
@6D(DZ5FZ\B3YR&ZKN]S')<&Q08EG!3E^)L_XEGZ F>T 
@XN\N(.P8X8OL?6QHK@%QJ4A>]KMM0L3AVG()4855PW< 
@?"2W$6]O?"^VM!P%:BD[1TM*Z.F+\[-J%'ZM?,6M0E0 
@ES_WF#Y4-1O?[=/K;^+U\WUKDH#D1/VL@YXI%557?$H 
@VR]?:1>&W_\:):H91I> B1-%J=([5\CI->-B$4)N76\ 
@[X)C,:!GQRT&7:QM@?B'U 8E!@0/@)7CAA1,V/N$=.T 
@#& S =I>),?*M_@NP> R6Q4D22& )5?[WY/1K[? GJ, 
@OX4H7AM&;"B;XG%/#X9-)LXJ+,9_ 7$AD2 ,QT@7@8L 
@,P=A7+UU.9)6&O-%^5ES8&X%NJ/IRDNQH\,B/ \4V9P 
@=4M1GT">OVB!N(9A/(Y7$#7."]L)I3:\IE@&G></2[< 
@S?F11T.P\%L=,8(LLJ[[*/I4T@36#&A)VDT:'Y#=OQ< 
@>@6CB4&,"#?0JXVRO<7"P %G3OL#E)O4NV '*O6N%[D 
@^]">@I_ZV#;4RV'W6Y\,:Y162QWP=P1&_D^ .>VNEL0 
@9"F ?$(;BM<UR:^W$]1I7M'\]W-9]VSI+#P\.YX-5?8 
@?9U#,40VF59&[4$",EBLOL,,:!#DS)1OM*,X7C(FP24 
@+L]T:]]UK,%,(6[3VL]F6[XBNHNC$#9_T9F?][QU$*( 
@O*N8?13L%WQHM$ZE0Z7N8C""9C+M*V,5]$<Q23L38.L 
@@,_\U,C*JOXP^\&Y0TH(C-N,\*GH6Z#WJ5B1[T7I=8@ 
@NX4IB2%OV\-6T ^?571N2F&,^YE,=1KD2=@B_TAE5!8 
@*L*U@E!,T-L%=K2%"NEZ.*_LJ.:M+$C3S4-W'GHH?_P 
@^A",+[VEH@PSR\C^$HK^^%W4 =*AZ]RE>7;W#?#^.LH 
@[R9 *)K#.'7<._<'/,]U-\2%95%MNG__B=E9@(4Q0,\ 
@ ^%5]SIR&[7O9:NRT#"^2O")\D6R7*K\SI7.IM8_]2P 
@-1;ISARD4S_L0YON^WXZ<E*+PS=^RY/S[":)7SJE>#D 
@C^G"K7YMKVCHIW=3U O__$#:"@><K'&CF.U</&,#5#D 
@N3>:MR%'8I#DQ^[#;FUJ$7EW54 ':_P,Z<&:7&P[D5P 
@#*5>>GN#-+;JKX418$-XX=3I(MD77 >-/9>&O\M0X%D 
@4(0TD5#?%VZPW7GW-Z,YN5H@723,$*ADVF72$LAF\Y4 
@O=Y/BL]P_5\PI",:$=_#S,^KLTGG$,;.%-^Y UN>D(  
@W- 6\]\ROWL-7M'<U4\OPFK:7B6K$BAR 1Q;T09@E/( 
@1)9.URL$A@0R4"A)4X@?+H6'@"UN/(@.ZEBQ'<[LG*$ 
@@IA@<;8'NXEU%X-T74*ZV.<5 6R ?E[1^7>(EF)-(#@ 
@+<B.[<+2J2 RAQ+]R]"H<O('[,)>""C;\3(?;0R*LSH 
@Z+G2'^2DEZ..$ZFDJ4YTNJ*$=<#;>(NF(^GLZR&L,)$ 
@<>21?(*6B!F9T;Y^BI)+&S5$C3FS?NA.6*$R:'%3_@X 
@Y\T,Y;$Q6*;".*K$R(?.A))P9S&"L=^;;HM=?J;$JF( 
@K5)4!H"H8'[NW'6L90S6R_?PMPM*K_;)-QJEE[HVKR  
@[.>:CO0N5C\/^%V/+OLIGQ ZGSON N?LW9U,,4JAL @ 
@]UB:S]G,421&4U0(OT<40?4<\M?+@5R]+"OC('@=Q0( 
@4;BS66_\_M>P1B>AU]X/<<1#VW?7R3)FL%' ZT[I,#P 
@F9;[@ANNFR1O]W_A4^6'=%Q]AW/.)5[,E72"XR7W.UP 
@%5" R4X5W4-KLE8M#0W"&PO9^7T.-,T9(,W9Q1H-5&8 
@??1BRZ[A@2G,^IC5$47AQG&94QFZP?$ZQB8[=&D697D 
@)YGB@"PNA4D'[4C)4( +5+<NMQ2$2\"_>OPI?@&S^P\ 
@!I?3\/PQ3.+.F=5@4O-2/UFP)SLCD3!MZ'PN-")'-+, 
@+35K[,CJ02/2R"F$.1I+<#N#.F#?ICREUY[*4[(@%Z@ 
@B:_03 +(,YJVL[#5,/^:@XNL/V=GA3!YL >@,7?5KZ@ 
@41IF"\J\]X.<(.%9V#>2!'9'T=+S:"_B4^X#\!'ED;D 
@G%*HCJ\I&&HD4L-Y;B &P\1C7J(4_'K&@MJR5E'8_,D 
@B6W-3.V"V',2%]65AR&,5S64BTA1\P(1&8>/$7=19"L 
@C_HOE<K?:U"+(%GF!CB/A*BE5_M=56S20F-WJ(16@SH 
@(8QY%Z[$&8HRC725'!G?D:/9J3%L<A!VM&YT%G?YG$\ 
@/3>>R%(/G0Z@2RG_)TE6:GD&Q5ENL#-]J,W%\X?=P?P 
@#1X7,5DCTT?[ANF!L(2Q,=,J?MSRN.<XQ,&?R@<(-DX 
@/I6F4]W?GT*?;FN@2R0\^DM_S1T(IY#),W=DAI=7\LH 
@IUU\@4SQ&<9G#-\%HXO5Y,I+P)R^.=SK6W[>;[3U.^0 
@VVK$?>)V?>9R3 KF%M<.5^3E]UEU&CHYUO8T3_D#G&H 
@[FM,>1EM<+LNS[K#9CS$-C OXLF ';)5T(H$,P6KJ@, 
@5%337'K%L%<CX@70/0V;'3:2PW_C9:'D'6JE<$VEA=@ 
@L?6/SD4^6^LI!2$68E!2]C%TL<E-$+NNV5IX-NHH*5( 
@#$D4U@],8IV$=4D?-<\!,,*U<3^COV=C33-[1T@U3D8 
@ +6;4>"SB> D>^-%&3QY$B8"'F /\\+1P-W#_5<0-FT 
@_\W\$ 47^ K)+.AAY&ENIJD6(C27C*LU@'8/80VCGF@ 
@E_*AFPH@D98>9=P5ZVV&$KPT).%AA/Y$8B2</?OZODX 
@W0Z4U2GTH'L? UP1_YQ8X2U]/J1IY"6%NVDGJE[5G@H 
@)A@_BW7A4:AC,I8AWZ AN3R29W?I"$&WNG_#P'O2*B8 
@H]".6/IDD1CO&T$BHL1:!"FM%W<+2_/%-U-?&:>F #X 
@3; _@( JEG$%D'KBJL V#42K A@_'1I2SK;LG1T /VP 
@6B 5+Q7/94ZE"* U.@6QF<XU0X\)B/_MMGDS)WB:J;8 
@.!50M7ZN])2->5VQ,8%_SR5+ C][:A,:'9>Q\KY<>9L 
@1'[&%GHG5<(9+T@AJL""9PL<#<]=?_6E):U_I@>;KS@ 
@MFDY2)%,F#X/.N>VM#CM;#X_BSA$M8,M+^U1O)M.$IL 
@$<;QEV+=]+IC7[IQ7%I^?R:A?_0_0_*(&S?RP5$]F.0 
@9J;\?DG6X7G%!'WU,TH:KA.0:Z_G^R3>A63%V!$II[0 
@6D#B!IX:$5T94=R=NI.0_1FC \=4,]<V4%/!/@+#_K  
@!H J6:.)..4 ^?456[<W*7FQQ?IS,Q\[L-V#GGX*5UH 
@QJ[MM^*+?T$ =QU5QARA5&KCPUSY[*J;*R3A;TH)L8P 
@:7)JC]"I570^G*)YQ*CZ&#G]2SM,"62G\E$\ A/8IZ$ 
@_O74VA,";T>#W>R&C8%C0Z/Y8W'MD^QM*'67=?C8J,, 
@K()Q+YSF:F71&"65*P$I0:27K>>Z(0?&X_>J/B7?_C8 
@-BG9XXU[N4!R/@OX,93M^"KT\@7%R;FP0T^<O?YB-], 
@,NXEYNCS1 J$'KUH-L.DO_;!!:4J6,$Y'+8H[ZB]XH( 
@J2["AM30L!N0V,C[WO6"I[4HY^30AJ; A.=<5U>"1U0 
@U6P1_L'^^TSO\'$V728">:.TO'R6]>"'0U.?6MZE?=, 
@&JNX95)DQ[9%E<X:RE9.JZV;0216=\-&++=&_ D2^K@ 
@BQ6[,]':F[V'JM0FZ$8CYVKB+$T#SL7[E"4]6C/Q>*L 
@IK13.RRP>)N\E"J*;C\$EN:QAO=UO(GS72)/CXC::0T 
@OD"5Z9O".^Y8:CV%('4@?@L,GB0+.3CYQ3[FPEA/K*, 
@6#H8$Y5\-R.RY-RH_)> 'VW5V%@+MD$5EAZL[6KQEO$ 
@JR:Z31^@#/'"A*IAH%$D>C;K')Q;&U\QUQ@!3BO][O@ 
@@KF>U<+&91++&_TRU+!;K\&@J(L\_P:<>D06E4JOH"L 
@"2@S*?>&Z5/8XU:$(0X(61CGS_T#[=3]#/;CCH-Z\?X 
@N^HI_ K55RT7TX8XB:M,V=SQ[:-/ .H&_XG!2.2W#0T 
@UV@QTF$A<*,M>.,^FXFXYI68".HV!%/>J#42-Q\3R>, 
@%!JZ@7,YQ3U-'N"DIR[!JY*6/\X/QHQZ*68>*<2I*J, 
@ )- R7 *Z2BE/OJJ&BCDDT'=*+-IBTS[H*#L*>-S:EP 
@[T%WX30X[D#$+I]_^$S"O5X#0XA9>7:D+;EX8?QH:1P 
@/E/[:W16@*_QW*XHYKK//D^[,;5P=RO%.S- 8E=%*BD 
@Z8>VXCI3W?VQFH-<L_X0!K8L>:3[_@FTFK>EI/S6,+4 
@"SK1%Y;XZ*W^4^D\8Q.GY3<ZMO8K-/L1N9^@;#_"'X8 
@Y-H<;X)X^T[=<UG$P361*X-8,*'OV$[MNQU& *9;QW0 
@T;G@N )DR@AQNTQ$2T2 X,4_65NN_U9_JZV99%WC)Z8 
@W%_+L\DK&5^?1 B+!RG_\]DJK@2-6XV;+SMWX\(EI!  
@ST2];)^5WR(-JBMK!-RIS[>C7]F^V,,!JHP\D+!MJ@4 
@MU[T0Z;"*]GBT)66?YF5. PGI'$M7=M$8DD":\);MZ4 
@,!P%\E40>WJ5$+X%PG+CT82EPBP1H$1[LRU: ^-TEPP 
@.>U\GV[K@DQIL&FSI'F#,?3_"@&W?V\SW8)*/MG^F)0 
@%V@#'F9@\^E+:!W!,:U$44"PU43-/AIU/W<^<KR"C/T 
@YW81O1VFI?N,_DV<Y,+E)4_KO.K9S<#&5Z/,PJ57AV0 
@*4NFT@\SXXKY&(H;YO-\BYT<QB_R[HW..\-"J;0=&ND 
@$)%,@,#2N':K>)+^188I"H7*FZ[M<;(,RTK8_%W"#%P 
@\.'JTK);Z+Y7B8N<7&//SDFW;8E!T8@B[/RX'-44T>H 
@A8^--O)C4K)KU?--;?-S!4C<^@B<?Q',R%-(+%?AK)< 
@=QC[HS"'I"YMA85LK+.C^.Z6]';X,.R $^4@4!"Y/N\ 
@". 3.V(NWVFI[>??;J'!"T#J)_Y;$F!)#J^=47]&(#D 
@AN$L+G%Y2AN .4Y-NE?Y5X&4:D+ (W7Y#[)9"V81S^@ 
@3J2LDI%^#]X=^T:);@B0;-@]W=M5T?6?K0:J6H9RFI0 
@.PE$4F_(>^C,/DX]JEI&JU>"BB+-%37G"P 20EAA"Q8 
@@S"G+:!KG0/!Y'/HX^[>ZJ^"T.NMR'?(DX&J/.^2%ED 
@B ;U$0<X%AB(EF;YTAI%/\;$H<DG*<9^0^99[49T;_8 
@W'[?O;36X;SP:FXB\Z)\!O76^8V FR;1X,)7RBV5SEH 
@BBT)X@2RB5M56G06@,>_*4.<J?>A>,B@!C<1B:W?E@, 
@PC+IWQBOX^MN$\9KI27WVMCM[DA<[26P7-S[XVIX@LT 
@SA.M;>E3_Q1VX>B;7)WT\$J"5.Z7NQYK&%V.Y!BKG)4 
@N(*2_1A L 0M5$< Z90WG6U\]Q7=7:=H91WW1B%\0<$ 
@;I*3H&26^^YJW-'$FMQ(IWW+A8M0!*G1Z#4%74<$-F@ 
@BFJ.TG]>:.TFKB:\^)-69#</U<@(^U:LT8OZ1V;^\W( 
@1([E,'AK%WYC,>P[HF2G83 ]/_<;&Q1C83I"83YB?QL 
@0]6,5S;3.1,7XPFG#2#[JV(Y)$1A]\*FS.&:-TFM?2, 
@L"X9U.\>*(0O-CXHP*JG=Y$.PC,CW$T'C<A_?X=-7'  
@-B*388YJ)7 "T[XBF"G%%63#4_O*L)43NBR]^O)F=F$ 
@%AA$>! A#?<,D- &LP4_1IMR(ZCC!W6^S"3_<N*4(JH 
@ST[6U>B)9'+G:4+88:1#U9N7;5@49S-<[7.XY4]T;.H 
@8LY:=C?!C -:/H.)7E!KO(58&$RP<.F]+$R&B=,1V;, 
@6GWI,Y;^<]Y,IPOXUR$K06)I70(HE4GMH$ -M2J4/$< 
@^E%5;G3_E6.GEITOK;ZKA)#<1-&)6(9"EMFDM$#:)S8 
@<C190T!YN3;#<+!U(N"D&Q'D$.T>U%B<R*UZ?? IT9T 
@]&5SY HC13PCY^ #:!!H5'1Y,Z@\^Y,Q8*<\H<(#9V< 
@C/&<NPV?[=X&+<8YYXW5EQQ;T"LZ/^90#UE"A;QE$E, 
@&,9]7N#+=A3#]<KFFQ+(&GV$O0R,=NRWK8\?P-^.O/H 
@7IXJR,;03<B;=\Q!%_##HY!PV,!.AW:$>%3R5'O^P%  
@4:;@5Z)[ .44-HD#$%YK, %(N,]T&))6@N^ G'Z(>_$ 
0$+O1Y.<(H1O)CVB8*?#CU@  
`pragma protect end_protected
