-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
ypsYvn7wzNP6/j1gKzMbyyhX6ZPETTEDUEWgS4OtH/PL288DMdKqrXqvLah4aUD4
B/n1bOq//AvJiGSkfgw1/ymSCnI+8igEFRkH65d/UD//oCXp6aPQXTEDsdRgRMkS
5Ke1Xgo1duKIhKjIYYxOmYaI/RLiKbPVsxq+50gbDALfIUswvmlEDg==
--pragma protect end_key_block
--pragma protect digest_block
Ut5C+3vyD8haKLR9GLesbzKo86I=
--pragma protect end_digest_block
--pragma protect data_block
M1rM1U8lXjUcu4KobcHIeRWT1mBoT48WaL2M+XqBwUaGf9fxfHeCBwO8Pz3TqOZA
1h0NVlDzh3JAE5ENL1VEOeJ8xJ+OImHoDmyokgCN15pTYLyOnWjxO8MSh7uc3HGf
sGaTlaiynYwgtqejd8jdHVA14mqA72XC+BG3BFwvLR1tZ/YB+SCc4RfKa5QO4GLr
Hq768m8oTQn/QrO46iqb6/MOe/H1E3MRKJ0AlzfWS0qIDFH2/FxJlObzGO85I2K7
TTH/NemCbf90wB1igXHBF8LZdvSaufSwaQI1HdhRbqQ7Ty90LgI9KVwE41fx1xCb
DZIny/RbbGNt1o9INAkgK+MInrVaDhVJ4VSHrmadNu9LB0QXcW1mzUvSUJLs/61n
qhH9KyRfjEzX0zEbk+a2i0YJCCjJBumyRyDyPCv8lvSO++S4DsvooDSu/DdprW0A
xiFlDkb1I8b0PPfn5T6BQUpZ59SjZq7jpoOjaF51JMJxPjagpUzWulIxGRIhShY3
pt1x5dYAAHMmd6vHKVesP5p56vk0j0HGwHzn99TW/CjK6DcIW3rrz9rNVAcvbj/D
504MmZY2cBg+wjX2yjikrt8fhL+/eKaFMX8SxTyBpBaCxSNre9Hj1fFz8fYAyEWQ
TjmrgbdfxFgZn1CAuihQ4jmzXV1B5USwJa9ewcKv7ZCBsqcrP8MT4pxu23kGWert
6646tF+7aFL8naaaUtpYyy3MGLDAGc0S0LWoqpwbNiNi4p/NlU3YLrORyHgvv4jC
Dbrf90U+rho6c+dbUqy+NtoYirOjTUIaWYglUjYRNPxElpD5kLck2WMqiXaTHkLm
7TsvWF7r637BaNNxLvoXjgblQW3An+k23r66FeMMBFteON56MTkbe0HKuInXexSc
0waCgkOHi/c67RHDRK9VzKahdBuBrXHE09YiYyMPGG7p6y86v+XyAm16Wjq+ale3
ql/cRzXAA4k0TVRU8sEcL4tHYZd1WFysfUdwoA3lJF+g9oHnqDqvSieeGNS+Ep9B
gaJZxElN/ql6D630h3VuK4/z6Kd+X0DghSgeivx6CulGIueEID754kFjT+aYb3jA
+JV5urGAoS0ixptZFB+xfPbqzkhN6jKE74ISf537ndOaMjpqqge7/oRzYw4+ahMc
CK4ds+s1zsOJgMpJ0I1cd5k9ph2nGJx33v367jNEMk7tuFL97xC617aQPlFYUE33
VVYGTo/C+u0+Vqg9hIB5Z1idN5Rwq2mKn6zpPjkgKHEzfcXD9ZbOqDvSp7hU7cqm
sXdQvci9bOhY/pY/dYlRO2TynYc6aY0xU0+SczGgsIBC/kGqN1cApuuEKI7ewNff
7V15EKhRgHKZ6mbhvos/35LLJwdHW6HtMhYEFSpN20gumZDEvfgiUIdsSCVkwQDk
xtFH8qg1eZfPIHl6KzwcoGGrN5Y6SozUBr6c0tSg7Hz07PHHrHpU+nqjLYSo86p2
fh3F9qIUieg0/xOce5Sy+l1QvcEviJquP+sDAKG+gyEgs2MXGSbhS3IGtC9vfzco
x6DZ7h88JHYHhCCfF09CVUyRFosMabXtDur2xUrorLbftCtW640kSrA/+bQ2O3bd
LKIumEKpx7uW2q5jyfzWEakkW5AI5KRFUBdXfgB0JXuDt77wyNGFRTPtcgzg4Got
d7IIfdL3M3MvsQ+BgM7BEJAvzlg6R3dUdWWe0AksTJ9xA8HG+4xQskPQH8d1sez8
MF2LA4Aivm3xVsePr04YvXo4TtqzLFH4K3YihYzvc5pxaa+znO6YhsT6j6UHX14x
xiXbHMu6aD+xJfbkKecPtqkmmrjTFfGTAmCOtWuAGkW3HMxbASijpysPalegdSUl
jaEXNqCLtlvECmxo8Y9/xyAYzVlma8gSOfB+kbqbL+Of6hQMcgvgzsH4Y1dpzEYD
lvA0isazuEP6vPjHBzApzzR+iPLk+o1zdiKA+uh60QIpQuFBI1P1I/CS6xNNmo5J
tTBOdv/49fOYT+Vc/Zhy2XXcK5NrZom1SB5qMGt/DnycPQ02cAExgK2+H96DGSyp
s1Lb5PI2lRaL3UC0nz6nmOSMjEba2hWBua0jjX33f9Tmj4DiiLtkPdB2vzATVFTj
nAbeh7m55f2zAOOTLrjBmYdIUZ1Zq1s6SdR6iKH06PsGL9do/smbtzx3jgfuedlJ
kRHPZbpco8Gsvj49y9d30u6VlZe8FrS0KSn7frC4rnh1X2797NBppVRYzUBAgmcb
BTQNuJgzYWgmG44i1xFckPue812/2GuzzJCVSE3jq9LfcUVzCGnGxPd+FamfgDFs
BrWHhBgzY9hP/QIXRGGYcOvS7Dwex7W/4E7xY3Ya4KjH+hcdXS7oIhjwYo7p2Coa
We0OMFoBMfpJYG5K0sxOHgnMQjKDmC/ytam4XXR+gtDzSD9VEj5p85XzgSVZvi9z
Ab4jFhOW//JH1Haex4oCxEC6BmQR3q1NU9BVjbDRS+BC2FU8zjHbwda4VQ7SkgUb
kRV/iYeXkQmdG+ZbhP2BLgk6uxt2VmEgaBWJR4GUejH7RJZYQu1Lgt5si8MBDlhJ
jJg/QqlHr41m4KYmVxZjAyqoP5Tq3PiVlAXrLWbOaHvH+XpoqzUBbCYLqBNt1rtZ
vCDOl5f21EsrzzKdVB360F425nhb/kJrKvR5YpAwKclRmrFNTc0JXp1abkOZy3tZ
qYoswyp+AL2GfZwoTUQSoGR/wgBubUzHYbAQsO6YAw1Y6wvxxwC+M9X1EjCeIGNQ
STatxW/PwZOFjODl4FfLHt2Q564iyK7602WqXRXf4EvMqK/y3CSOoNl39zHEDeiw
9vXTBHk6cWb2SaTWebrxtNoBXSnEy4jVCA14gIS9BOsmUfzI5mxD7Kdqk9wDxKRG
UJdgAqQaFPBWU4PPisig/O0KWVcp+rE73XHiKR9XKlGNeGQjw0CEUM7Oito8mVxR
OZGaiR+z9K0Hm5XQ6marOBPM8ixQeQBYnzDWefl99iylryDVOWTHn7EjQbbntp5l
4oyTSrt5noraGZwhWLQAjvX6+FIxhk0V8GGOPca6gxE5X/aA0YGNCgWGrOQPsjwE
1g63z9oSeAmpQCZrjkI2QmMQvPm8obCl6W4U+I5HqCATxTG1zSmI2n3RSq8VmxIX
Ig5QntoxLEDs5CbXwq/pThSgsvMrmUweauhwjC8tY6Z+wYwelYwn3a4lcWALM7Y2
P7jmh7NfZybKgEvWkwJ2tkYaE6ipDbE/bY1vNyTlfanzXqqz5KvtpIBJpp2GQV6S
V7nxbO8KMei4OIiR+1sHlOttncniot3KjWTVxfDW/QWZ9D/aeKNAcQfiLPLZL+p5
FAOXZec2831rTfofGKwlgRVm6c9Au/F3zshNWCjAi/7B5EPRIurkcSZkM23ODZbK
bly/bNrkOlaPazBhSFLPFD2as0FxzE7Sq1pF62gacV96a8K+w3lsYH3J0lCUJrmq
Z8PDTrQq8U0t4neZvCo4xetDwJr9F3oINsAHluPGo7phkPIO/k4JfGb3l0C1pPNn
cgweCwzM/8y+B7yyW3A/xRDwTnxnFMQtm2dahHtTQr2FwHqSfX4WWF6Qvkdz5E+l
HVCi5sMA45gwf2MngI0XD9HwgMoLj0Wgi6JJx+xln/DNi7hWzo6SDPD0oalHk7ra
fvx9aVjZVC/QXrFbknztbEBrwLEpY752TWnAwmULxmHfN5Ng6zf3X281b9FlFbH3
6EbViqmqvsTZ8BZjIyQekBi04Y5N9/tE6Vuqkcp7xKjJwosl+T6c0WSYhoHobmN5
0Bfls9KW3QkWJF84c4vKKbeXNEGS/BK/1k5atOGZXBtsTBdJq9jnozh36gAAsApK
UESLwBQO3QAPyHEtYQfxmJ7k0wJB+s4OZLu1lrrcL5mJnnNu1O8tQ1oz/XtbnH2b
I6SjXXxMTN5PXf6FCphlNF+JBj1gjqLQz9stZ14Y/plNIz5etEEyWZZqYVaYXham
ZAOT4AxhIwecdrMNko2CzbqUwvGfaKKu1lIJXAB0sXSwQ9vZqCqd6Og13wzra8ok
VvdyiU6GLQ/6Y9Q/QMzEKWlCVVKovHBoL3A5PdzsxgslLQJ7lM1tItDx+DLdyWAb
kBbnf/XwZb8Avu+n9ucvugXtIxGSvxQC+Pl4XN47q8+F1aDkyNMzkqZ1IEjxUSFS
PI04ammlSvc8SOEFuN4LpydnRFIzvrRzDaxBFiniP6O3BAMJQ2+y0YuJDjFtwOX1
NekmL6SMhYRCzXP/3dC7hhAdicXArw+/fBWNd9FqI4Nru6MZbKCuHxr4mbqdbIqQ
84eZRkvvM5eF2OgILk80C3q2oYWNW/l42pp5DCPhYYYKkGuA4bdQolm0hQboz5tV
+/16CTYLABoObHCFHg2m/pMUZRgEK8OGEe4hoxAie1loopyLQz4kGTDqvTq7CCg1
r2MoT6IsmYNytLCnvpBZBfgtcviOsCVlkyIQ7ojqc7QXC+yAH1JLQPxoBMEyEhOa
WQOtTutyRfc9EthkrsipRBAWPzF7gcIUgCxk8NsU29SEruJDEVTzqCtbRLJDeWC8
cw+6w/aHS7pc0m/v/dpv6Eoc9z/LSEYH0oyWPPRdW0m06uK3p2oSIk32PCykKKGp
D6AgTRYjdk/irZIdnUz2jKJhV0j9EQlIftdLbYZf7QiLysfBwbTCE/nHjd034PAn
L1WS1/fAfwMeeQ1jRRZLF/0mSE8eY0+65jIbY/yKitrMvYMciudyMl1YCgqZ+08p
IfAEJnIsdFkuL2M+5bLjwTKhcQ+o6bxB+O2mSYHAH83Ivxq7tBBcDgmURDqAARoU
KiTTmucRxE4khHdMuFaQ3w6R9/J0vyU9BHEwyimldEsMvKA3k69oKa58fIc2H71R
omtbT9X/kNjVedv0wQ46vmn3Pr33WTPkxfVlH+jo0L+AbyfOLvNxIskqMNl8uk2l
Nag5005qy3I9REAEPwYNx18mnP0pDdRIFw77Dthu/OBvS1jKvINFsL29VpxPCRWw
qKvxgVGeefLM4GlKvCYDTCp6/gRATPet3WeyoNfpQ54yYE3MtwjetUgJAC2bKtjw
Mntr4Q3UqIxDkI79DV2AV7faew3QX+bCtVB0fXm/f2CWBKTMPWcZk8anj0aU7tNa
B83EMU9GHn9S+qTjxU07Uj2u+s1eLFL8KD1CeqSoAhNVRkKRIGAt3oE2xZn6Y5HI
wslRNIMuGOjTzPxcycfPRa9fwkzAs+QcVCTMXCmzmX5tMCVEutTLE5Hi4W+7PzWR
8HVN2er38Io4UJzbfgB2PxMqdGitLEvrleCfxVaNsv8cgy5vv3UN8oQESGpEvYig
dBfkdoV+RQzviXxZoZIdTzgoktFQnRQt44xsOf03K/W5LVuvh96xnektozv23WLX
6LN9arKubOmJ6deUztjn1DvL3Sv0YStlTIF9hhO6EOxJk4Yxr5ALCmJTLzo4AQbP
TuqPFVAggoO7n3S8osiIDQyA3DiPd1UVxIppvfVR5vq2V4Ny6v6Wfboa7GfgatGQ
aMmJIpDxrLZ8n3De4SgT40VKTPLSe9nqTA0CwGBczQAasuOFNM4IjkZ48fRc9u/H
bKX3Kl0PhpWwFesilf+aWUYx2JUVGsHQ5vpev+SDlkl3c9YGgFOsFIg+9s08kIwt
BtvcK0rkAW34p8fNdACqUjykUIUGZ/m3BaM5pULy1QAD0+VhygXJkuxsDpVPo3XI
stlKOA5zOsZey73zccxuwBkoAlfsGZNTqDB1FHsqcxByKU9XugtDCWOlGJj+0mY5
9JElBa5zMn1hPXdNBRMKgwnbY4s+PyjhWEdrDi9JOEaI67qzbs+SqenYCFxevxKZ
Nc7bxrGoEAIFe/Usy55mKcrWzNtPzYHhgIALrJlqCPWp9i0bESHLL7Tfri3fs3uj
9cr4ihhykkyB18PisNXFikasUXz7ZWLckHAC2foDt7lQw/xN8RXq60gVR81b+aPS
Gn3nDpPnyaZlwwtjFo9EGSyM3ttUsfgbJ0U4dD2OMWZB9f+GX/Z3CewQ8XJEqqK9
GNXQFOsLE342Eh7Y7H5PLlu1DadqIiPLwR5cz+ufG1C1PvA5SRaJfjf266jFWen9
D4VlD1DJDvaw28VS6qM9p6+jVIIEjZVFy3BkTLnwBIYVPama0S1vhlGbMiXShYvS
GDuVURDiArZxHiBBrv1/+vLLDHDCAzgpZM7vnSjduCprjlB710guAL/p5g+yN4w7
kO6JGHbFo+ycAwTzQATTd2IwclMWX9WE9BGAp9qzasC3lE0VruFLPFlcZQ71bvBu
Ohm3qKsOeR41Bvqf/oO6SV+kAWeGmtJSDUKf6qUzuSDmbYyXj1AxY5n2E8AnDYPv
axQpFbM4o+Hyp4K7/Q4artT5VomaLUmegOILm8L5kTV8mWcfGN+grNPmZhg4Zt/3
7+GZLskcA4JQTz+9aeaKQAtEjop6wv50Yefr2cWlbWpZpZG3BdlfGMqrDaI2sOM2
hUe+QvvX9yCFD3j/1Bg2M3KFUXc38CtrgExEsKUGaiIjpxZ7J9Ws1SMXPuDoRGe3
aSJW+0G9AFP9EkkteU5N8RuuMIAEaz1u8Xw8XbS83nSUOg/mt7kQHW2CB1eB5XZD
aPvnJs48AhVrihQ6f5E8rPWjq9x4skmcpWxrvSm7uQNl5Q9f0NPcfCGWZHwV7Znz
YCoZ4kak0+jUkMdfEgdS/PfJzXaUkTJnzo9r5cL8Fb95/Q0gsm/2vbiQuoyQvJsD
1ifAxuKEz5moB/LujS7lXQcI3TXUzgXs46WMNaVEiiNpBUmVdnvMZ0PRhVcWCxSf
KZ6lN5Y13lc77U5PrH03N01009vRrKH0/Qg9Dk4m86E1pP1DBhiCFceR/Pz4+5SE
Aae/pMNZWKGdhVADfxj/OizrMpI0m125JRlFeehImGuJkgsnNd9WGNzeYvIHTGLz
U0nd8yZTjfR53us4oWTagCPM8LjHRVYwkh+Fp8E/xAkzMMPr3WcSMXEbik73CSHc
Or3zo7IdTySQCifMHDyWki6jjVIMoR6cQN3i+8BuXpA5SzOqYZ0Cwj3eVgI61Mdl
CCoPYN3P6dGMTm9E9XtoZ4+tgLxm1FIb9whDshFkJdnW1P5uH9SL2vXLaFYHY5oW
Q3LDc/HBd1F27oMUfpHgb/wg6DqU9c2DK5OkXtlEyt9BSmScAQ09bJAvMiMg+EfU
vCRaScmsjnew54DwNa7zLk9k8hUp9paoccoPfwp0RWbGia0UtDnfKBlFT/sA4AMq
xyAOmsSugH7gh/7tU3INdkVumSJPO9imIUN7IDlmPJ+mvFpLXxUgX0aS3TcjkfLN
omiVmCubtIEqGNHAQ6gO9N5/r3Anb5YrdEjJLKkU4MdX/YyHh3lELUmPTy8PbJOy
mamGTaxzqVeRSslX333rLoz3pDGCB7pH/gEeAGx5UdEpJktGuDetjHmNnwJXdaMx
A+znIee1z0WSm26PcFwKVV+vdVSVXZEDAPgeXnwX4OhXUhnTr+gWz6trjZ9cLgYm
mCKwA2vqPVcaf1KOj+zSdcWRynif/BAkSMA0NbxMpJKdeRNdvooTAGE6jUC+afGD
K5z4umhQQiF2H9oBAUb4Oi1/eReKIpqnJCMT/v2eEerYEgy0RjDWjM6kD5NN/EX6
utnm6zHsXZFtWiR5vSfMVWXa7X+ntE2h8nuiTRoFafKhfcdO3T+NKfEbeFMWa5JQ
o4R6NoZdclhQcfmrJijCRSIaWQm/3FMJ9NRKvlQyji/CpD3z+kmVRmqlIaHgqy1G
ain4gzuSO2SzVGYJkhvdUZNu9XxCg7IT8suDu6LuF6lc0CxbAN3YxsvOXVI8A+Hv
qZmmY61yG1tJomb3+LFrbIOSVPRCxWEXBHsN9wgLFYmp3l8JdHgdH3+h8bZO6nAK
pECF5NBT8NQkM9SAVskatp0g7zCjPRwuX1PRSMhB3mZN1MWhyTPHeKOwqQQ7UC/K
AYqzw6DHYhHOoHyiLa0n+uGTy7OX9RBa6WhJf1YUetJI/109nL1KyKtm9NVJsoxW
DpxqhG4XiKou9uPNBldq6qfrBnJcccjaNS3H2q3ipUbMST2TGIm2Q85PaaCoi7c4
4QbhIL6M3f5IRCbUJrvvVeaRfGNqU2TAhMm8pX20TliXMw/GR1b3rOzur7nMQYiE
JX26XuqTG3uAbHAVB23C9qMY0uCVDtoLra6dehFu8QaANtghokP6FcpmKb3a6Wm2
32KcWcR9mg4ABfoz1Ktk5fzRAWTSA0ugFO9dVebBFfeKRVHcaYLJMGrh+hi8xe8t
q/OKJg/UCXPKlVbFHEh94byUU3haCFLrmZlCw/ysYnpu7/9Pmy4bhjANgZnLlZJX
QrRcBJe+7krzSKCMM9+AtbcXPn4mhOrsN2MbYCjX30aSxJyb9KfmayBI5nFQ5ZR+
sQfUoRAxSld4rHPAVz2MBlePMDXslocqLKphQih3Bmqv1c/k8A9vE9p9fp+I6+dG
g/6GNTGr7qsOtkZiHNVMfwbccSQ6tYulfMo8Cpg950OYzIpmIX92EZZhdIXbsXtl
vQIs/KkU+6+qANySgMvuQxbKao+6rfJ/W03I1icWjp6hmaEFzyyhwntJFypO92rr
M5BS2Qd2GzfQLUfND8bnC3P4Wu8ZqdV8CP/oW79kbSJhcWrjmpusDfBVXPU2dF/q
dcTi/DyUQSEb4TzPKrR/q6vvz6vvEHd9wCZLL3ae7cAxdKEQcySC5wVGfBGMSCkp
IIB4LeXteHI9E31OK7oTnSS8vhDosL9k2cJmw2U2VlZl/O7CMpYJkCBmZxlLsBCp
iArQ651RohJ+D90nkz8dNmQ5C0AqEJH+essd9E9cSegIXd3hHfpSLOcrj6Sfbs4h
opm1iim0H5fQtjCZVg+RnUvEoAkmISJONMb6RiA0QXLXee0ik1e2peDw6Rqxd+IT
wAZMoCpePLszB4KPxuYwOruXakAkzVafF8vX+lL7QYmC/Frn3sCqRhDLKWPcHas6
v/t6hLtmisYLQGMG3bIZlYMo8MwGJvGLbs7H/ZXEukeZAy1eTPVF/vBHC17fUXe0
9t8OHWW+4dZ3Oasd6LpjUeSb7xsZf/zm4KLMUp1WstrTkzx49z36Jwf5FY/UOIGl
jgvFJ11PsEqTGHlVUEXyMsdxjlYxxL8LtcW5t+yUs1JvTVt6f3vxVwpsh40jYlOV
GmQ69rR4JFWefLpPqyLzhgkrXTsHZm94e+RRlbnycRT9ZcxZJe7UGxGj+Tux+kHL
MXHO0Zcqi/GjzPMJDaZrSS3nFdqwpDg3URm5g/hl22oFdvcKOQCIQQ7WaDhvigXc
ZNUgKDCvi8V3m8CMi+JKOcccSpHJdfUzefnybbbwxbDeCNhRsbJQDXmT8A/BrWo4
Wd5AeX4YM/1mwBA1vUOe6A3woYAuosgC2xrHo19o9b8aRrgiQPPiwSkGNuN01A8h
8/CP7vx1RjvRSNzENY5W38w8UuSS41XUE1fLolOG3gvoWAdg9B2BWBiTahqsSBz5
aHfOgfLFkJwd5XjUQrC9Lut+j8Su9tyPFdKVoTnoMYm98lE7gq7FRYFQktN3tlo4
kPJikzibaU4JRUUcSpYjha/XGedGI3a/pgcHNfgyzNZfof49Upo8eWTFPWzNKRhp
uyls0G1IPzkb/M5xmwOutWgyoqa5vDlIxWVQw427cZcOSZ1PKn591/wyxpS1kkCq
CjnPgEeR0mYWr52tbxqLUTh5+sdWQscx4XITROtjfSggJyw6ceWwRjSxW0hWFad0
rOPS1EyGCHpr5oCKX5fRzgInWfv6L7uBTbSHHfCDKctY4OwHYfTHUBcunFVVtTtO
+jRfk8F9zwldnoOnr6yqhcW9F4lCdJOlxzf/wHs6tMNmnV8D4VnhWUsSQ/vR+iZe
WI4IIrjN+DC91tYwS81u1mLQbbhd4VQI9v+zuuN5Dbk/mnftuYhfxbUPU1kak852
R1QkDlFyiiWhC1rYIlcXr1KFVhTS1xA+sLQcZVFh7LjswTI+mdavQAzboBi9bVmy
VembxrvCXSsawutInt8QK8Qfirm+njMIuy3fTSASVD2Ip3EigyfFtYuRE3BxYkOC
pGzoC71X/GtIOt1OmTvV5D7qRc7uL6vlm7/fotoQ7bvfU5K+RttNFwVoJd4xAOz6
CNK0IyxkyyctNhhKtx3iLEiDaReh+WzV2aRb2IoXM7/NuZoktxQ4NNrsyMTfgrKY
KsNz0/DZ3sQkP7IS9jxBTcwWV2yPGsNN/+0wMbUc17q0nBXoBS6XPDVCrZiX4YhP
2CH/mZr+X5y8VIZQ8inj1IB5JFo1s5PGwXox5oNXYu4=
--pragma protect end_data_block
--pragma protect digest_block
LbrUubxjZhsNYbjizGsHgj2TC00=
--pragma protect end_digest_block
--pragma protect end_protected
