-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
kq9qvA7eZfa+oyTWMhCmwki+hjXEingBxbBPHJ6BPxdd8ECISOue4/3w7mmhLpPx
E9F1LnQ7n13O8x4l+NN0WY4xLJ7AMzHSy636RmypBdkKfNsnyfApCugEzfPtKnfM
7iiGO2KvSpvoR3TM82Q1smMtF/TNHfjzEJNmM0sRkU0JoY+vXHDyPA==
--pragma protect end_key_block
--pragma protect digest_block
SRx2j1N8FeE4rnMIl/Gw1Lqb57o=
--pragma protect end_digest_block
--pragma protect data_block
A+IEDMYLoRyl8p7++8oBp2H6Wuk4NW/0jEpdKzC07xyl1aP9O/jdMcsT8UcyIN3u
e7T8VpXk55PJQ+xGQea6rA4PLGI6mbLd3+6TAk61voM3wPRTgYdsIDnQjV4AQhW+
BZg86QY5ZS1WRQ1w3pdYVh0P2rVUb5sfRNo1D5u1dupBy4TxZRa+I1jjTAFKNeWD
6K1Ewc+Eb/lKklU/RFD2A9OqWjgh/BGequf2rx5PJtU3PggWfAMRZY5SRXGpHvfC
5jpSR++0q6RyosEeBTDVfgrvRy+0zxYwDg/fTJTPPjfC8j2+AfClq8CKdhbN5q0F
bM/8xApBgDm+dyLyNMDMHiZNe6c/w2ewl32YvKTu4ZP2DcTDXF5mbJIDqxPFUff5
2Of5g0N5PXbAtUapAS4y9Sn1/Gcw4X1nP1ITIbAIiLPVouSyZRG23iHpeX6557k6
rD/UJdahiZABIZ7Do5UQNku3Q8sKm3iUg3JPvUGTN+uAd6T3SAePuh6VyYmdyUvg
4XvbIYccXo7ZfoPcQI8usH6CvH+WITTuQKQ3dmEssFqEKHdSa3pBTr7eGO2LFZxG
Lm3NnhR+IjecGxDVsAsWp4EQVrrA7lQONzhTBRV3egd2cBlyEZOWpHOIO6PKVXli
YbZsJ3vkPLH+Ey35Zv1FbdHjXrcsQt2k5GjMaZW2Ya3oppI9U4QnHVDsuCJL8pGF
7e/rGNMOqdeEIygzaet7uh6a5cKbt8q/XG64Muu1tUuMgFxM9lo3emSwJk1/ybQI
rqRqsvG8a7VEyfAGFoK88R7eKhQShft2eF8HCzLmCVWapOWPhaAB25jSy/3W/TKX
s2tCgPzUrmk6xBta83FHVj0bm9k9BVtEP5KNgjQwutstbKgOhV/YHXYRo5yxRp2v
CFXaFXR4akR/cSPP0nWZvDV3Ucuw62mrznWCCtzG7pSzbmH4yu88uSSDqUQWXSFj
OjixIYsQmTPy2HRv5UyKVYYqJIpTOK9lvpAb44bGkyd3Ylz5mQ5yHWE65MT++IQH
BLqX+SPscUtVvcxFn2ofbh/syvtrehsJ/V85M6ddf7ORRE0ZsL1fpxUpItu7xbQ6
R/0PKulRfXpUuAT/WE4QyIBBtHX7sipZu1CF1Y2w1DWVi2HFUIJT93AydGA9O7Vy
YmMosGxS1wTN06s4nOedy+vt51T0T1wzhAfgVHYMTwiGO0yvV3qaSQPv5zBXniT9
/iXpnZPsv2NcPs+gTMchAeNGD1W5Rf4xiYof5oH8w7oqgO3CaHiTTbuN990V+ali
gUVZsk31igvcw0uH0wV0C3y21INi5a8nHiOKvI6sQaLSrv1wHfwO1BNhuBEf8n7U
XiDZlyW7X2XmuVnLdT33KGugC6sNDzXZKUYj8VdOTuW3G7qbk9UipBkolDpQLMTv
ag6r/yWDBBZEbFrVeDLi2sVMRjX4xIBkZvAh6wfm6bNS9lCq0sR2+pXw1YxRjxly
WS8auLQai24/L6po/AjpbBLtslt28xKh/XGnloU1qPgsA10c1DbDPrYAqVdFP0Ee
59BxTazAJ2ROn3EEEncD+DmMN5lMD6qAOzFkL5WNz4wZacN8xWO8baysrDFhNJiY
zpSj1Ps6ssRde5y4M+r1J6i8611wNZy2dabFEN7rhAgbWBhmiIA5rulwXkZ9AWqi
HVxBR/lElNDKc1/gbJ4G1WalW9nXsTV9ZhlIizMYIwu3e01F5NCuRWYST7+AMQjF
gVcYvWZpkNxiKcZ9n81fE3x3uFpgD7qEDk4/q9yOhsEZsdjj4qBwCi3xGTnb6cXo
KjX8e0gLZld+9DZhQrQ1pw7FpjP1sFIH+QwQwECoTVpq3OzekKYPqq68NMuv9Feh
7B+EEktH+KbRDPAgjjLk8vhLtWF6koU17ULqKfO/aN3luCw/Wu1lo9WTBzztwqxJ
UEvloNzW84OAMtm2O9PkiQLUX9VVIF7XUuxn4g/CRPuil3IAyUK8gaBHcaiGQUGM
WLO0WKoH3icX0uimV1CRHcIW/OEHRjY6U3byBQJKO7k5emOP3aH6Clu1BxUmYFhP
D9N+yPzQtnNJTtHhsUCE115A2uo3kx9OCLLhUuAVUEyYYYrBoLYgrfI/ElsrFYdN
R0ZX1FtL5JV0q2QflgP3vRSwrx3ndI0o5TfX5w/ppTC0XaeWUR2dEZSwrUsqNaOU
3BaU8yTPWWlnDmWP8s7kdkHIr5k2PfD8yaaE96zoYjfPymRGIenuYv3syYyQsiDW
n0hmo+6aM+H7QanxNQMgVtDeSy06h1Fgd9EsoeCcvGN0XGFwcdNXtve9v4KxjM/B
LjNmEvMBiPCzC1hYWhdrTr2ZHrCK+6QC2bJKDE5mwdssWuytgigFKOUaKdMzzZ4K
ng2sR5KBGmFeYmUHnFO2PQerph4ML+zK1tVnnX4jOL6bex9invXYfU6q01zs0GsL
PdIqroBNZOwDlI5WZv5h7UEeMpIVTcxi2Y3SMVP2sCGsLFBoOquh4wM8x9edsCkm
W19eZ6TD0q6idKSv1qsRQEXHAG6NHA9I5dlHPyZn2jGYOtYDTD8b2cIiHE8apGp8
6JtukD/37sVRTmSc8ICWWtk9eFftuVBlw5ACXNEWLI1PHAwg/GIU1XuRA/urWEu9
2lRNpAN3AtHBMpQRE+Rbmx6eW57dXuBS/vIGEq7j5PUMSf/CAxKechdNxvAbai02
MaD1HwBTNd79s+/+D/FnbW8gWYMLnxxsZ3AZWc/1AcRiwOan878WIhfCJ4FaYN6C
XdR1sNiHymBhwhD17ty+2UiWjwGrRu32GM/IEhLypaM+N9Udb0HqkHefKslZJLar
QDZPBgThryraggjCAdv2WbITuqG8N+DucGPxIX7KAa7LgAmdq0JWVXUje/Eo1b2m
I7r0EjyYxE6oj7fOmIFr+s3RqUO/G64vmYvN+WZLI9MUTTve0AVehLmOQF+IxJsL
YevMkx/FQE8ib3OSMaiTMUrlL5kbvyL48W95ep38vP/E98v/75MwLgAE8232c4JI
MhVA3NhQZf2sJIn4byhIy0NULVw2OFAzKw2yqpILSbD7eOfbTEtqQaD+Bg3eQ7M4
r2u4YqXVKrmQHX1IOq/OjZgHB/TBQasla5o628avU3aFTdFmvpiQx1qFnARUfxHf
4Ke8+EZjXuQmM7H4p5GmhSHB+vGsPlIlgVmnYu1LtohESSf4pxGJTjLtFTs1ITjg
P5PmyZ3E8ms0xnH2c4rCROAT0OL9hz78tuRqFGhsVVsMKh2YjrFD8QgvnOoLlQVz
KI3WRynR7l0E1Qo0KYje5/7Si5MHQ61IEFmU8wCF4APG4E/cLomgLBpLPMnSZB+F
b3f7SmqbZXczbNJPv2qxzpMJcwNbxPChFh9dZeW3D5Et0p3lV/tJPXijXg2edNQj
Ce1si/Afic7JmupysG2V/Z33MjWsnbMqSLbGVLq1zQXSC7nmmVK5qKjjqhWC5L1O
uOaQZcGxWv/xPNNgPTfLSG7TarSVt5OhU6uthWzJ9QNJIBFq+fCfbwICGnUzjztp
RRtZQ/vRMlMVNAhBTTxY+ElvfYwrtJTSOIfWuxVWI9rxLxmX3l2duMg7vJ8tyV+R
wEwDmmxklQ393z1c5fk5ltOEU9ISi2l8yLk0w2wUbLcxa8Sri3NqDYTxkvhwinHj
atV4KOfCyJ1oTMy9QmaVwL/qPEZhI4y83NLHyjJsf0sJNHYjl21WFA8bWjXTua4z
Hnq1h/L7upggSoC79fe9Ohvxq1R8pR6XuE7zqK8c1v4keLUJnO6yrx5/7GRb9X5m
LMdZFmlhd0962cvkNuoY6RfdiHUN+Fv2MvKUU5nZtw6wWIlSs9GFJL18s6JZBMvI
ySedynm+BS6UKaFyV+uBctd+Z0xnUjfJHXXSKMxtgejZnroqzy/cCX0YF2Ey0c3j
SNTMIuL0iSUN67STgfUj/JMXhVEKfaOZ6UlA3NKHUWqDHRC8SotPWo8kLJQeWDDA
Bdu9T6zNrbFBtpHBfE1xKBhGdcqbr3Qwzb7TK1ft7xGr6j6qEZLjYB5ldED7QGBm
26kBlJzcnS8mX2nP1WiXnQ7DrvcqV1K8RYLzzwhu5dW95JqM96Tn2zX9eW5Mz59W
vFMiuA1wPBjZ8iwn2/pOYjkzzClGiuIMNiMODgVEry2/7wpTpdL2ZzeQJemDR88v
lCFPb6XX1rbwYtYX19qeYmHe426xePo65vh0lQiQrc5+FVrcqfFwyLRrBVB4HkUU
LXx5a1gxupDYs3leaSAD324duwbwAq77L5O3GR+Sah0zjdha/Hawi3yTloJDzJIv
hvWK6fP9zlts6JfYnHZB2JKOHZdpmbjqriWCmPn0ozkNuQNOWbmvBB3tfheuHsNU
YoMkVcLT5NfrOX3fcOMvFOI61dkQshkyCp+V8Hx8pW54Gv6SQ2tUcJ/DhZG9BOPQ
v0nHTz2TJJ2llLVmZjGHuGgknjpLtPifxian5QPW1AtcOO8bklf5NW3YvPKdgG72
9jSNrRDQLsZNsBzrmblSYzOCxGf/izwmfiJKEisFa/000MkPFjTYa7zSoLx545vb
sOTz2Rj0k8X3Q6rGhvHB7Ces5hbq1KIchyYCbxX72HiKFTIkSeuOnmK1Oe6TnnZ8
Pc6ur9UnD9BEhgSg0tWzp1LNW32OiYhkKzPhZ0cncQDfva2D61svaE4NXB4KfVY6
AndDKn6bL3OtE/2fIbvLtwoyUCx6xab9YAHHhubJ4WHA8AtWhU4POFI2puXhgSVA
FhwMvcOWlNvBZuBXroQG5h145Bzorjs4/anls31zOfiPlcpVmxQZVDgivkV3Dr3F
vF4eBOBiMWazpVtr6+vIjGFop3dVGyXxDJvYDIyFLTai2rH+lAyNrGXylrO4ikz5
tcizuqjj8kXOaIzgN27Wy7t/vPQmJQhtjvqA0wz1Ti6U+Z9qCMcLTC/pc8btZ1Rs
dx8dMv0vkUC+DRe1Aws61JXEbzIaT+c3q6AJyjSn6a7NGsXOSeEyLA72HajktfNV
ArrCTGrQB3eaitsm4p+GHx2fCdM7Go+KbQkx0mH54v2l+U/mRYGTUFMFvtHuagvQ
5fgLFwFDgDPHyA3uAMJL/rd/lGM4VtyMwMxw8iAh1VWaThn79/DC4bJDTWv+7GPT
fDGc1ZqaFBUVmu8K2b5UbB9fwcIhIywC8OtehSj2gi6J8ptzTu5dmKdDxiNtXDv1
x8n5PxrhkkuOxYHYIDVgkdj2o5Nt51pOk8NngVKDoUg7rsgw67YLX0kZOq5O2IZI
Oj6dE+M+DySEjvKRZiLLErCkCPyhl/Z+UvtWk8Dk0LLeEZqTf8GZZEVVVVwySTA/
ChEkTWe5RteDUWdg67Pf6ErFtceUjhnSuHtCQEmtD6Bp03XByGZJuqSKOWJdtgYO
dKxVKrte5dapWsVg4TDt9rtf2XJK6Q6vMl7VThHCSBRdO35oVVlbMX96uppSyoGE
ImLlm8HuxZX1tcF9HwMfySVULbAgVVreRYsVuWC8DEtZgfLC6EcXhyVBS0a/qjRX
txnOhbw1iizEmLGjpcW5TzeMeXjHUiNxpN3bgMsp9HJ82tN5LvT2/pS18y7/hk92
CKPjaCpyMXJroW9F2xnSWwSEmzzbsd2A4bDu/dO+/JJtX5/Dzr9LwaaTcldvRb5U
y8qiBtIvQicqy+XzmYD8ZRypfpHoKTeiwzYBZ8PFoZr119oPxpqBXOFKhUD3ZkV5
lFrfkRp1qc0LNx1xbrT3SXLTXKVhsUii68pdNQkc5c9CGFYk3Gkl+k3qtd3ET29D
jLWOLwKLZjuODKkN4F/zAGrjo8qdrNd6JEqRoyxfkpUKTfWffPgQwVDDsXGNNj+Y
QNzNPO8Vz4wEYBrogms3BuR/5UAkbOONqNq5AP2tciM+D8X5Cyp2kyg6ThWRvC7y
ldE3en1V9Kql8WWGJt5gfEhhwB2FnvWDWG42P/CMHyBHi9ITP20+qgIjLUJKH7E7
GrtlWJ0d72+dWwzHTcZvhInxVfMFvsL1euBiLIMuq7W+2/7xweis7971jtXNQdlz
jkHiWUFelNv+m60RSDDyALgd6l6nrHnzgekKsNRibRGayzDu+wUxlv2kHE3/lUzV
RN4kUoczhW/pDGRhPNqqdkjev1nMH/xRBd3DuoKoyy1uiAb4/0USDcYRIfNLuj8e
wMHWBNK7/mMLl++hnSgWWMNkNhd6YZENuy0zMERT70u1/rroS/mRbC2t6sptznOi
6LfC0aZaFLNYxH+r5oyjSONVAHG040EsW5eaFEQ50ZBmEyh7+mOHkcwhsovm5wzf
ws+9/YBJEG1B2KRcl+QeVhuSP4MLLzl5DlTpGEXeap7GgEftL54K9zTipqk6gcXL
D/5EEV1d01wmCiM4zzNYMMb0aALyREosdSyur+Old7QWdwFJWtExZ79PDHO/mnbA
SXLxUJyHK8zS/r0vZHG7PbOkOjqC+YYujZITbrAHdZ9bQpB52035RjrpV8A4N8cn
SXrZJehEAKzsGy1riCwltrZZRZfUdcCSUxt+OSkrTm8rfniMS79PesWK8VQyMvb3
xT2p5GNOgw1MxXO+laSBXaiXNx4YSGQKmMf+mhVPXsd5nlYzMZnCKEf2+uNAreiU
lg0b0YbnwV6i2CXJUKrVX9JRGKF8E9G6RUSbTGc/rfKKVlaignhe3JH7fq2cD9Ed
FGKKoByOgv0TmKlG6tllhg8v5WvqcBv6Mw2oXVHqW1u/LWkFeF5x2vMdzdQpcqe3
gRNlqoYoWdpw5fuDPOsr5xrGEeRVeQLRYDOHKZbtDAHEc2EGfMWCrZ9ARf8q7XzG
vaMlkMxUgZ3r3rANM4z23TNw/ZB3EUuhWwv3mP1GyjDjvB0DeB0LnfIAz9BLuzMY
k1rXjBmvWKP2loShhnWon6tEiv/sZ2ZJKq8NaJCo03E83PwlWeKs2k1UBDHqm24b
pkbvoeBd0gKswStC8vkHVJ+SM7hCIiczMZJQBhVQ3k6QFLYK7Z9cbCNGVw+NTPI4
GKi8+7RPrq2SJhBqW1TkQDnDs6D4UXZfTW2LtvvPpJSTguI+rrkhZ2iPPmUURAR/
3S9INg3lIXWfRfm/cYlCIeWZFrYlcQvr1hIgTDBZdeXM136yzJr03QifloCbGeii
iV+buAvKHwAkfJmt3gncLdQAMbN/CwZBAxNBOCy7QrgKW4+Djnqn1en0xcVwuJIw
WOsvsbRo6EB7G/Pf1hMZ/ZrdifEUaBZrmhRNWqtldVbYhS9eyfDavcfye58Ff9im
vnySe47L+ltL6C2jXXxKDpo5chH3Kp8KIDszxAgroMbT0VtBFjKqiTqhwhWwK+ph
gTGqXkGP8gU/vv4wswhyPXXylA9Zc749wqb5dT7xne/zxHz7AjsU/Nurq0x7t9VL
1Ozkeu4g6l+MIahFnGTzJXdTuYYLpiCr9QlUlQJNw4E4A0CB3qctk9zSV3+o5OHv
1qt8YIvZAn5oY6DqCHTocZO1GTUAUaPKgphmzfwxGPNWEfobTidW9RfiB0Eu4/Fj
Re/fxMAMa2ep7hRGHDxv/HEeozpiVdMDN1OLQgzSyQtysD2CC72CTFXf1ThgCX37
tHdNzuDA+odQqqHgksZ0Dk7pW4yRxWOIdoHQGKvHs86CrNrQA/iUInogMgqRn2h8
2t8VPnY9rfqXTXhQd1gCM/iLXZZoekJv0Ehu515LmScRPUKfvME6Gw9dDAF46/31
JKUlysOG6t0BekQ2k4o9sAK3Cpv4YBk5awtSzK5rIOFBrkjYo3I9e/2mBFYEZpxO
6ByD4JaPqwyo7vUdxP3iaTXeS21HBNN10xdBJ9h5Kp2MyGRSficfEHb7bb5e4ddl
xfjz2DfDhzJAI7sllmrPE9Xn1QwNLtu7MJvcAdR/WWONO5PPw1QISJETvBjjNBiF
Lv1OxNt7HZtXydR/UoRn3Ma2Vt9hf2LmHIHRMgxaAL/F0uQ0IpfKpDgOnKpKrPlf
/bdbOCOsb7vzIhYQuFxYQ91giCOljrGGyYxjsqhL2XJfiU86rFIpPRmOwOgbbRPD
B3EgVa8x+KQMn0j/LNk99gN16nzGY/8106MqHNFjLs2XB2roiH1lr8kpIOYZ1Fhq
55OjIq/ces+oih/jl0O/Tc/GPNOx0EdIZnpYe3N73i5fRm2cN61wYNQky8MSFLZb
6pg9FuBHxN7RHo8AbFk+ZxhKZ0iNxuMxDuaY8xuDLPQg2jjEFyotAZbEOJPMSrD3
KPEGDSLRkdTr1SoG1DVTtT1Wjj+Ayy1z7AYRLmOVkapRc4BqK8O78m3Ch8AIRj19
8iCf6zYPSaTGH92MV15RSwTbIw5UjG4MJsFhJYXCUJGDO+E3DifYnFM3FBAEZ/qL
gzC2Y3ok8m8yi16lqfmRhk3NaNFdQhawdBX+mEkN8vqp66M5t9GyaWt7u65CGq78
YBILLZN36aTzAqo2edue6B/ccDKZiiScqhx7v/yIMnl4AqipJ6dHUoa0WdSE2Jsy
sdUn620oGw6y9kgVowYFlmMG0s75X9+xvGaviOS9WMzDc71i3W5pZSmEGSJdMh/J
X1zER1oi1CkSz7m5STJZ2XdgUjkwQ2Rive925+LpbcQ9w1bJXz6y3xl1wvDyZSle
m7hZP4LHYcEETfGu29lT3KQJs1aj5uZBiex0cdtcNiTIgaL9lpb+8K5mJ0emZfCL
pZyaZ5g5vBR84fop5X2Z4kTEAgXl8FJndBm85Y2uA7ziLKHMEgJzRZODgp+5IOYm
cuBF+Ob1ARtirggTkdVtLRMuhAsnFx9h/IFEL3OUF38KUZqgV2O47BQCrtYpQzbB
SEzsTm/HUm749h8Qbu7sw0ETR7v5x4wWsmsNQGF15Ai11jbSqb7gMP5u2hHvW83K
OFqbocpj511d35K86J0dbL596JPKsyKs0uQEQaDWfBW5uD6NRV80DatEXxwsBI1z
sB6E26KSTyxLsRHs2vTJg2MxeW/2l/XX7I3K/kPNEtq5JgqDDUYKkMiznmAuuySi
vvxbN1q9VaLkIxbWfMh0zc0Pe8yYrJBl9cZ3Mcl/rq8tMP1M43n+TdahAjyijQKH
N5hgqlQ6NG0qnhjDWoBxUQFCcIq0Dw3TfGD5GEBsojCmtvWHymbI6xL2eYwz3Sum
dZqB2mFVCuNe9/E9WDeAUoAOnLfkBlzFi2U+rV+xZ8tu9NWXnmBlGD7yb/wmFKq3
Y3QHq9J6qu4pMnz1/aJBnez142hxZdbisnX59uVySoPKQxfOE7vwnae81oJvr285
qFSEJgsD2EIKZtLuIPJi9mlPeTYragOdbJTALAcl1EKqHzndcesYDurF1uKb0nWP
QuKknXnILLXSHq6CepXI5y4BkI6qegyAmbKP2pq0ouhcn2HWUdG4eTgJW0xhh6d3
W9MAC68cglhXci/HUEDSwu+fu8uxe1Cib4P81JRBss+eYYU5bwS44Xi8G34fPkdn
jH9HKX7pbRyXHRJUlICoppr22m0f1R8v7ISiI6KWITKjui+T72PWSBCD+Jc9z3vE
+F2T/psA2dpNOhV6skd5hfPEup8EHK2n0AXpFJjWUqoJuTGzKIBrhVCDXmVGPPGf
XUIaz6gPWDIFsIxLAgqjDph7Ch8BlXSyI7MlAjfpb8z5Kcx6m58xOWI7IU5K7hjQ
ekjfQtEBvEnvopARv6UAi0uvwY2iS5Ox5ISg5Dcypg4Cph0neANaeO4ksIeosiuz
XAsOrsVvZa11DD9iEbHn8DopKGuSwdHSyryBrVNKmCgWIQEwOQb4EOCkYjF+mpyx
cl5IiMYImKbctricBFMUo6vIAwoHwIU+Xg8s6q+ceVZcsUcM1RUF8l6hfA0IP3VZ
fSvTP7CcCJQ6wXAxBQtv/KZ4iTYlmRFMKarWva6xAYL3GvydH/GT8HfvNgE15AyX
yX4hXjwN/cR2llZe6egpXHhoEykvHHGdYeg0YWLsvityEXphrO19eWnmMDXiQy1p
/FVr5ZD5iDu6jqICkESnuNJHvTESCpZXxtVP1reAqCDm+e/q6CE9zJm7JfwNKrsu
RwB5SshPpvQX6xzhFc58XqzETlITAy94pPt2dPXWz+C7K9mWjnEtJaQdf5+6rYXg
YTiBsnRciZUep1UgalbUsC/UJ5jGZBsJVzziaPpONhpvorXbdwh9oL3dyQgx+2lv
41A3FpLY6G43OaUjTb3V4VR2tf9Yr7jOrNTmsr1DxI4aOf9Be+hxPagPPoS/h6zQ
tv1RT9VYo0v94OjtkSDAF340gmb+kojtBMCrNNhybsRZ+8+xSclDmp6w7ULqcqpa
jLZKka+An11dh+OmnN+2+1fhyL2H7GVrNor9pV1IzYpW5hOsmgadaEC6+hYozS9Y
cNi2Y6SHxXtK8iv8L+wsKycuzEdrTqOaAaPvkI39F2tgmtKR6bGbeqbq1/6v6UDh
y7oTAuUJEFQ+BjgvxMw1h8WS2lCwjJW506qNlkgpScColka5/BokTdU9ECfLLNrA
voOlYLRt6kLdaIeBa0Ev+aQyXHcs048uDw37IHUgfyzDgxyu3VDarSwPacNV5NKn
ro80WhcqL+Yq1dtUcqZ45WcoS4vPjG9P4VXlkvLsFYXTONvAHUhSEC6kGjse/GQy
+Jq4aLBnTh+Xt6PX9wrXhur23IeicqKFZGa87P/4pe5DbeF5t2spcCohwlYazPOa
JE+Ueg1tiWruVdB/ZcYsimNsh12QPApYRUY50lGcKsM8gmnAwq8lHlRfrxHHBzHT
iAtXsmN2i7JofS1hiH4k2LcDITQj10taPvKMnhV98yk=
--pragma protect end_data_block
--pragma protect digest_block
74ZqtN62DCF7Udr9XRaCyEq+EX0=
--pragma protect end_digest_block
--pragma protect end_protected
