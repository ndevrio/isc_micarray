-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
isFlEthTeSEsWNSe6fVIp5n1EohuEqkEwvmAG8TlF7KY0Iej/gLSOm4JI7qk7CN3
b1yEQhUsWYWN95NDFjniUBt3VL3xzxtkdsua7uW+cFtb/dxQ3/aE7F/glvbqEoSR
+0nieZVeQt6vAQO0ZlaA8jcRY9hG2KCTLjGMzOJ5Zw+2lXt44OIjRg==
--pragma protect end_key_block
--pragma protect digest_block
IuSTMXRiBAKbvKdAay4+/guy09Y=
--pragma protect end_digest_block
--pragma protect data_block
1MChpJhFVa10NCx4abWMaAsYTzwYgCsrspbfa9MxgO4y62LBJV2oVR1ZKMyZ97uQ
lIqi+mJPupd5/fRsNFsmj/+y2+3wc10/TP9fuPL7rHAyOheC6v6H5hRgc2acPnNs
hDIlSihY4si2bC36mTP4sSBQ9Vy8buzxnEezqrYgQlLqPn9+WLF3qHuRhVJMdA6B
OZOmz9Aany07t6w9+zB/2PkddG9MxTCsC85NOMI1UTKo/jTj3jElRUuWb7s6kTjm
xj/diyyqgDPxB3DWAOgvoS1PppBJCP7l2Qjj55JrIDAPZqGm8OQm9EYqpffCjPaK
vb9XkBWk30SKgmY6mVa25iSb2fgyDtgxJSk9EA7Sp7u4FIZbwjTAsZEgZjUYDIid
tuxXAKWfy61RviGIaBU9f6o6hLnGfUofAAyPwE/ZczUNB6uC1EmELpRrmn2kLHEt
bMM7nEE1k7mqpxLDUR5rGX7UVWZHY7K1c2CdlganbF77RdQMwAzuH2UaOxasRldv
zCJTnqgErX/KnESPVolWChK9HVuhUTqkvubqNX1QQP7eCwHefHZ/C7m8L6nDHWUU
hfitUOoDXZM9e1i4TEvbLSTiR39r5wVCAZfmnfA+VRQP6KwR18+mYlsn2dSpkLkk
kGTkGXWtYYiy0yHkdyWct8yg1DO58xxLmSBNOPszDvDiiI2lNXiiy5PCqh5IIZnb
lmOfiQqrfhlmgyEQnkZi9Qo9Mp+J6QeeHaLMGq+IrAxRZa4iqKIEtz738UtDsK4w
LUJNNDPku00WlvjcZ1vxmWjEWxOiZPG0/abtJLHmVFgpvaobVAD4lbY9T3MZlrl7
XvPR5W0nOEc2g+eD0G2D6kaWOBtuz56Yb/vhRw6PhqFj45zFoeoY5SPV66vB9oCk
51VVBthc+mi5EtlqEdarguckxX/tLz1wYqRVOeas8fGWufpuHiyTaDrw0rEzvzi2
voTraYefjQ7farCao7ex0eHOEJYPI+nhhTmPHf5mAho6JF912ThcHAGyPStYCL39
FtxVcaeXkn0Au/b6RPO+Am2xUB85Iga3JILs5bgNH6DB+oxKCp6ZAimFhf1sILVw
uk7+bb5BS6bq026PgB/2sMTFwksB2ZCJfONrAq38wQ+Onw/uzJnOF5bVSeNBqUEQ
Syx64QwC7mSrRG9K+d0ejFy9EgfXy7ejY1dg/0iRuHqjwsldjmtQKF3/yvQ4Yg6E
h1JEivXxhl4SrKtFr8uwgpEhBZ4xaNEmklfTmy4d3pwVTs2MS6QEmIlrGc7JFOxX
SAvL7JQfUNfniwVM6jzW2dHt7JXjLmxOxpTibxNlvOPbGA++aM3Fq/vCDDU/9E02
KxQusj3/CGiaUWZvYeIZXXRROje7UAp0woxR0jKVNHcN1MN56WVoSNfnJZLlROYk
QGaK5PL58/DD5jWTcXC6L0IHQ6wJFIyuRU15prbBgfRLQhEVlZbk+u+8LeBmuHLa
CxW3K32wQJujVJcRpb7dvREZCdn52j113arrf06/mCVLVBsOegXbAD96Ue/Yrw16
ZhxXYJmFuIKcInM9pOBWhb3Uvje4y5YYZoE7Q+izPucDOhbtjj2L2NbWPh3mQ6TR
e/Zt6FDyrIU3TD46rEQxdu/uotTrRaAVigulmEO+39mi+J1tAeFr44msrxlTSHAS
bBEhSB1DVMBGiXmTzoJaICsy3wTmrmBXL93lKeoPLGXq+z4Tyz4bI3o9yjlAhsAX
dxz43D4bB/Vp7HYVxMOmXBCDnclOp5VVc3Edz2crcL3W8DBSTMNZCd0bfVZ6tNgF
L1PFO5gU5fMnIyb7WPGU0VIJddPkO2gd7YMPdIctGajliaZ4my2HSJ6ydlRtXMyx
txvOHngT3KeNjcfoFtgoszP0To0fAxQrOlvm4tRNVB3mYHfxaoUgcsYxNCcrBUzW
ejgLnI0mKg0vp8eAELbHpp9ZY3/KL7Z63+L1q5tNmHH+1XrmKTgQTQNofnD+Ok1V
XQbyj2o6KaMfOTRU2wnqxWCT697cjfsxCaeoAwZBT7ov5d4yoRfou8zoExSoxLF6
JHTPNfTgoSBh2/FJ3Vce7ixfUvCbk1YCyDD/sZ5dXlxegHaRV8wvyNU+g+wZue3J
PWhmLTMSSmu0NT7rQ4pqeS7xbRapBvDZieotOSmVSMQggx3pThWXUHP7WsWVJAWM
fI7Wmj/9Yejwk46Iav2NcAEkjVDz4/PRn5mvn9K8aUz8yYx+xGA6n2B+s0HcAoq5
b6InU68DAFbzqjBOMwEBjqAKyikbNnecUptTvWaV109jSeLRlENYZk/nhLQvX1B+
Zf1RR9zHPXmfR3RYa+BPTI34MDq7NjjWAch4kKZhevJq/ZABuXmZ9i0oE18evMhe
6QEyIzhEelT8Mq2k3GkDbmmACI2exXplWQ1Gm/LuiVsz3mPmT4RyeYh4QU+WfOgL
qOwbHeRL2ogRielu29cUhc6B/SS38heHJk3wsinXgqWi0QI8sBVv7gQvwAYhNMEP
sOFjJpAIls7T/uFOcZiYr7a2Ts7/8np8i+3ix1x+rkX5cdviPYBJdkOSkJMywTEl
W2Eq/IyeCfAAue/ozVpvxA+yga4GOhqNArCsuJ1HI4/Lfqttd2Zv0pq2b8c1J62R
HfAbHvgZd5oySZjitWZ1XPz+PeRcEEa/suFh0STzY7Bj1/UK6f5Jb1uh0K3qqm9g
THWujCl48JqCGiPS8mGyCdtX5zn1WTGt5GxNJUh1GrrybVXZcAcPVDYusDkQHsY0
XoTvLrzJnLCcLkSacjvNR7MN3zUM9+jthgTU6Ol+OM0Quf5wld9dqZWyWcQk8OCN
GaRqcsAY2mqfUpvjS9fDqstWWMcgspdqKrm/dqYYhdapf+DnUmgfxrtpAJmyoEtw
0o4hdXBcIn+kzxYDwz5p4lEHhot1i1byGqrxUlYwH3cED7/UxsTuE+8Uq9Ue2Qjb
vFghHEGLv7ju5h+WsbsQD/s1wMqmW7fCdoLlSRByyZ7K1vhqmDEB+GQSzPEPVbqX
yMFRpXX7gqizTmaFVFEiuopKt6wf36xOsvGt2EIwXxxVv/ium8G63k7HhyfMy1nM
gvsqca9AZWRoC6vOQm4aJWn1rGYUXEmlbPS+JhszbD+abEVYCztCOBbK/Z5dTwsc
BUZdQERRJmN5T9Tcit+4w0+/2HUyqTEWCHuL1FZpYhOSTAO1JliZeRl1xKNuOwMG
wst1PWHLrfzycv/SOeArI9HrFx6mT3CQxwl9kPu0I3dT3iVT7RfcRl8e5kk2Z+0T
kNpdHNN0aq8zMvDjVGpVj5j4PNOSjAItG3GXVXidtMvetcPjy/AO0ez5A908C6A7
UQ8/XxiURJWHVZEHU1OMJTgpjYBZ9amylaFylrF3xc3ihDn66JrT1lBhf57yXN12
9B+LqWUGPUNHs60xj4fgw4VN7ikYEG/EWtmwvZ9mw/8u+Vb7erichplAs+jbqR1Y
gER/nXInozCXjiRKOjTiKCQKFXu+DinP7OhN7e9+36WldLgz/ZO+/XbQfF0culzg
/O2Ex6CERCvrhQrhAGuexs8q3l4TOVWOQBpp2ivAykwDayK3XDHpKMzPROWEoo/a
iyCFZLW65OiHO+R1gRYJXfgz9GuWqIesUi+/D9QAxv4yfx2laauFcYtKkU0s3WIO
lkmbDGSfy+O664JXhZ6vqPQpNbRt1GXG6+Sq1MLycBcssokeRnnwvzWfr2VDCc95
LDrMK4fqfaAjrVCkfLO8Miwe0eJKQ4CYbW9/LmikzM4OqqJggVgRp1bunwmKYeUw
fQNJy0uFXbR7WyeCemlroj5t1A+86P3ahD6CF8gJG11QY2qqp31CwCd9pKDsiESA
PE5K9g8Ko6HY5g8ghmOTQDK7PmfF7oII+mFQ56mOP0sUOR2Zimqa6oYDnUAW9Zkl
DjVA9QvM3p6qeDZJRHGwOQOgkqlrcKt/z+hA4uVVX39wb9TBRazJ2Lm1oGWqRmcV
n7DO7BFugRiatCw+pXkSMR39N/VD0SNf3Xhl6q66AzvD5IQ3xuIbI8IUXnWaNXzG
HT8PjmDg/6pr+nuRbf1XLroocLaWVtswcoZEgqITKWe3CPuDcF455QMK/0o581xa
irpwvS2c1LZiNpjWKmvV3iib0uHkwODQqpQBUNKweFpuvwkxjZVQ5uz+RcEVN6Qc
BeTeEqtJ4OSisOSxqsVrPSmNQyV5s+kUFmojgckEY4nwCzjrI3/59nbjEZjxcWlW
Xb4UcHcFiDAE9vCd1zjrWdvCOkVHhGi0eYXdDHt5+xsXOBfVqcOsp1FcNCpBpPm4
qvYpM+n+Dl+GacWuTSxBhQDeEmVaHekIJ+1unjyKhPIch0Rq2wZ7L1SYrwT9YO2V
zH9Uwf5CqpkXl1Bw6+iV6+3OSyUfs+NhYzqIm5TMeHzRABe/BJ3A5p1uEPS6AYtG
BHZTCkIDmn+JpQK7+oRFV9/hGplO8c0MJQWSVF6+cLfdqMwyKTBHngIWrBiMI69n
fRFRLAZeZsMeFfc24hwNBUW9Zxoc8MG/a3S2ypZnv6Xjm5Dn4Z2URoxjKxMM8sE2
+AlPAOdIevJy0M17/TZCdASbIknMUyZ8IG96wG2qFlaoqxcOB9UKOfqjImhGh2o0
P0CZ1EIECyTwHQz0vcjOG/dYCPXo8pCurwvItkfMI/xKMjFTy4g3qvG41v+8QKSC
RR+0hoQ/nFGXqyGOAJtONy45pm5hsBUKXXzMP+muwJ2Xihg0NOl1yGyxGtNC8WO5
OaEq5zSK/ZL2GCFmoegptq5dlp89T9HYMvnaBpnP4Qmf7y9GWi2tPeCUgl1V/Oyk
Gvp0qBOn9zFskX2qeGHHn6fJrCBRuOHQUcE8rvSo4kiq0VWoJ97pq2mzuNJJOh0N
kxRjZ+v+HPhs4ierl5Dt00rCHz+cuR64mAfmeWBv3WOaX0CI0sXZ98MZEL+qbD1J
ekQYGDANBeLFDqu4qzJtAvPlg5+tWZqwwoElOQ23hmqJxVbMm+QGxOFPyQ7s2svh
1A+qJPKpwQ+EEFgiu8xHeRLpCjWiEtz3zJz6thD4mGJWYH1Dmrje9RC8+0ZiSQiQ
xd+mBlLmVS3SGxLmaSilnqhk0c+ghYJ6+lpRvVNYNreUxLc9OipJTbDepbal31lw
FGnjkOx8w7MaL9/J8L/5Q0ojDwpEtbBkZRF4m/u9BCvYevumrWMdwaABFbxN3Vg8
GitXCgkaUfOR24WSh2g8N92tkQ0CFDpFa1X48qf9eOTeNA8XeQNL2DcBLHRKc75f
/UryY3nwxOfkePXn6mCEHXVfPcJyrHGSxDEcwva90UuKXg4JNE5leRE9oPO3vG/4
P80O2l5dqBra58NhWhlCXXJgXALsfEgiIFdk9aFEqrc2z2rZcxIoYuL3m878kZSA
vaIX2JnrgLH2rVGcZGYSrWMbDhEqEt1tjcvzRr468IyLxqwd59Y0egqI2UoetT/q
lLYa9qCE9zHkW8i8aulxzyBTNdArmZhslQPufVS1hOwY4kH2YyTADarwmuRSiiOt
jHEpzb8Nd6dduLadwaxEmOSD7111NMNu/Ci8NgXQKTIJ2u5xUSzofQ5RVOwHY2CD
TLX8zov64rv1+6a/rwNYMZ7YmUYOdm0loj/pdlPcqq1sG7J1tcEwyrN+3b8Pq7Gd
bz3Q28LoSFzoLAtuD62s0t6AvircAm1BxiHCj+cOsIQVO78f+hzxM7si+EXNgT8Y
Mc9ITBf1aoEZuWy8kiY0fqxcwj78EzPmy6g1vSCZEYiLL7t/fIxPSERunUMDtS8G
Zl53+4TxSeIa75qEB7M3QwoYQKjRNgaA6KLPXgBRkoKhw896wQGKzicIaGCjZz+3
i04dunWe6zwD1XC/jB/79XAyFCeIGBtArS820fvqb7dPN4bFXIhxS5poqslvL8RM
MsS7WXLLK9N2eg3G9hW45sGD7nt5ahEbIjhGJEGQjaAwWRSqlz6UChz6pHlZ09Wu
M9dRI1KVkHmfly9YDK+6zfxIkcQEdVE7YpydTSWXK8RukoCi8s+QQEYMybRwB8Vw
oXYqwvpdRuBxv3zJ7QfshrvA1S6SaLCjBOt8xfIngxoGmct1kRrDOUciXNbozXBi
IyGvQEh3xyo/iJaNo6NZCvQoh7rM1ha5u9Q44WbMTTuI63SpI7VelEbfN5YVAgkM
nasB/jS4rCoc3qslQazchnrjmRBeOiejab6K6IiGcb0M9YW0y+PkTHmsYJIzvOUJ
buU3t3o3Ewa5l7nO59gbeANj2kC8rqpeQ/mDhni/eGO04vN1hiQyIga4i3mBGRjS
Fl0Ea2Hf+uSQTvgUhh5fMVeiiDJCDOM6bkPmvfKpV6iJfFCPrkvo0icbP2n1U7VQ
+m593JoUw5pmN4hMzMuVxq43GuSNT1KNZ8/NkOhblsH13YUn6nQcUYCpG1Wl09T2
Gq5XmV+19t10f3VVwtwyA5I81NqJKVZMbGAtSoli3aGrJBzu2U7YJ7MUmDCRX3SD
Dz80y+49oNVRLxVFVgCV9pnq2+XjbuL571L3Wo5HbnXyNhRrhhZ6SaihJ2A/AS2V
AM2ApTr+zQVEJl94lu14nsrZI+HNaKsFm+f9iEnXo4dc6ap1yVuEDwi39b8LdCp4
UNn2dn4tehNpXPy2AzhqbmX6Ld73AybeSKjHWIrt3HaFQ+PQ4XdT5eRvIGIjXB55
yleuZjJt3ns3z1iQUOo82Dq8y822+Z8LVc4Wx8q1/ziwje/zcVA5srqZaarCOTPq
U9jTbI7CE1wSq30LBHyFwkaFovOwvOvCH3EWSIIR1h1jUn2WXo5+d+B+ABtf1hQX
O0M1/Q/Sjr4KqKs6mKsEZfiWc0kasj+/bmPDlTwxDWrPYVhMEgxnATJ00Xt/VKsk
o4PtAQft8PqFjomlBwvuYYYW6I+nxQoVsuHTECoH7TXMDIIL02NN2OTjfpSkDR5O
0udCwULfw4fHgk8nbciNLisbgIVeyxMKOI9wfPqC1z8+YrnxSislBMZAxv+8zdl3
UV3I9LF6G5A802bnv/OkMIzSniMa8e6/w2Gh6ARzS15RDCPsCs3wT3B5aCH6h0IC
XzED4O0oG3AVP74iYiQDuiEsKPEZV0vDkAHpAzBPfRJDhLrZzU/mcPBJU2YznNeI
PUmJ7ZSiStlRx5eICMEvOy+QN5BY2xYEHOqNDPtBBnCfCOCGsVDXukQX86ov9WTH
uFiEzttyDgokKYMrAwyleVz8JTLnuOVJr7rNmP4MV5zb6UHTlUq5cCssp+2jtXK2
0o8DTnV61v/soP5cgxjBII45Q/m/JVbEe6zYDxJHO1XY7QC+SXtcyil0S/ZlJD37
JTqA6mbs/PT8zNKMZS3vWhXJqJCQRp+L5PQ4PD8ON/sL4Z/TR3cvbYR40NEE/nQ+
tKW8fmbD6T5EyTyIvoj+NAb02SU63AaFzM6imdEdRcAJx/QQDAqTQ94KvxMw0nC/
Dmf7OKw6QpD1ovjW1E6HYn7SwqXsj/B7+I3T0ogGElFFfWzUmtZA1SU0rztBGO8p
dBfetzWBs+dy+aUn+DUHj6cEw/jwaO9tJURjUEw/DTM5uqaGmMWG5X8sP4B4tcsz
jwf3l2pqC4IehKH8LtYaB3lUEZ62cEKZLrYXGuwaJ6ZL4PpIpyahoaUpl59tMPB+
P5FBVUU//qIlkCbz9CdZRNQoDzwRjrZBnSHoUhnuMC4V6ium4f20WfjN2tv7wLB/
mTdL0lH1UVT/vKQ2MpN56yJ2YnZOxHCxtzdhgidcJK16ExIddcHC+m7Ym8zEShHp
MNIuyrZKAFhBTAd3dTpSGe+jK+586BFw9O31PlnqxQeoBVeXOcUHKLjajXlsbJM0
jaR4IsZmrTXfGynTsMH8xT9wDJ5XsWcwfx+6fiMSL03hwo4bOxCSVe7g2FAWrDKd
2xEfO9Bj1SeHAxoJYLK7Vly21ByzLqPYDECvXD5JGFxjVXiWv+OekB4RMGlR0fLd
lCqbnV5WvD0h64GjkfohldXX565yl7DTDIr1FDk2wCz384ckVzMNKpvltiBDl5Mw
INR2PZ/wcI6WJ0QtL2D5PSmBFDHKhS0pJ9Bpb+kZ61tpzkHL5yblS3by0psYVpTX
MPzllpOb9+l3xAVPKECIdf/pZ+iKGND/UcJs/hy8qF92CXSjy+uvytt5UJIx341T
kAPwFEXJwjHsrhuxUqpXHdcdRQNVRCpX4LhepEEvkkAyif1XPHi5nwxa6it3kQbc
XzMQRBUtoAbqp2aGvpkNq52225cWSz2QgBGEKLxY9hepS6F598zxUlXMkh6+RuPt
GWZv35YM42aHsTsx/6Q8ZTX8GzXqMrxb/ZHdKZ9n+7tzodUC2Kfm4thY3kZDJ9+V
qHSI36QXr3ogjuSgfSwz/tyfxqW4RmIbBkatprP0Nn8NkER1Cpzn5AGmGXsSrtka
JNsNetdyu4E+MTEAW3ppg5Ms8hp979CTi1viSu6IDOT/nlCnoQhHe1lhLAOQU7lH
URLTFc/RirCOmrfwVKEZAZXAPL8XAPXfv0kO/CKfMzxjfR/eslURduI4Go0OPZr3
/Fn98ZYbneF7PUCGfid19MrJZAqAmFGeIlb6GkY1hQS4nSPJy0hwBAKFQ6HpeGa1
MgHNGSbLRotuZjMHeBd7992RQ1qF3Is4FmK6K5GbbTtPD19YzJN/b9/PyZT/TA1J
sDBwZ/LCo6NXUtjT7PHVDz75C0fwXZ0R9TMXcefuCBhYAyyqZhH8cxaxFYaiD1mL
0UTjDBKz70rSGEZDFVI3BfBccGxox0cMaZ0ZdlSJSvBmxh9zbvJRDUpW/jeMjr86
TNfE70f0DHq6SouheUoK31cKiOBPfykE0wsqSw6KfLzWaO122eXZRcePoFuOYdqH
FuVsi2mkmv6Zdu4aj34yw6NaksBSRP99QJ561mctbfUJWHonXBvllUnWRoMFAY69
VWi5/6Wnwhc7oVVZN6Mgao9N0crhGaInV/eCwVY0GwtpN/wsGUjS6KiAINCSIq1s
6iDGogethQwJS5xvsGlpHpAONdwvGpJQ1CMeAztnT7NSkULPFqV1Tyxr0SDrZzfy
eNX4VEFtsHDLDNsAdGOEvjtXHJran/EGx9CuyB5rAqKkHokJqMES59Rh1wyB/civ
cqLDWXdsEpV05Pn4E9hM2BqLpNHN/+ZCa6iEl1X58XLbBCOVBYOBBt9n39oOmQXY
aMNI5/TspRqsA3rfVXQh5cTZgngCVIw35eZDJXbx7jimAahxDpVvZLs6HJMR1hoW
RnDyTepkCpGOrTzHyyk1tluzGXctd+yepjTpHfpiVDViRYswAs0928rX7eBHKItd
SCKwogvNkWpgRaghqpYbR/11LVYHZnPCXSblDnvyZGfae4Yh0+TIgo0bu68N9WDR
D0FONLgecr/Pk2Khw+sZWjZradwtvGHRFNW4wZRIfjpfqlmQG22eEK2AWBOIBrP/
EPOvuIOjoL6X1gCgItUQ5asXVJ1FLZTo+gcyadBGH4zsRdUNnS6NeGIGN4s16H4s
rvEdCdKNYpiuM3eBFT5yAoR+X1o3hj6j7U/oFY54CWrOJ1GAheKOpgxVmRgEb/ij
S4Bg2vZBsB5NqsVTU3kyh2VTP6jw9t6qoIGNQKJadaRV790LJK8G5Jh+RbtPu6gD
/4cOrLWSsVZM5hyiU66hcWpiiROz00OWMBu5SPq4Xt28q9G//PPi8gzlx5E/QOSv
UwmkOi4QtPMFO6P/BFqc7eJurIyV4nnbYslNKCAJCl5MHv5cShfy031rrUl/435z
S0zB2N/M6G4IsK7JyC7d90MuE6lovmdIDc0lhuvO7q1oC0e5OY8bfFVVa4+pmY4a
FFmMrmV8gbplIaRQxtP6rCEFQdhGg031wdbHMj+/TylwPgliQycM5aA9Wj6V48m/
UIs3xs/9NJ/wvonk7F+LSEqt+5LnNWUVku71FlmVJIJ0iDMxVMesgvz/C4b4VZkc
jRbE41i4TxKqf5xh1I8V0B9eZgtNwQqFzTl0OKkWHP2ovUZG2psJRxR55Z00BENM
9CGJ1t7BEjTOji53MgF5FHFB3WAwtqZ22c4+MTYl4oPbcADw7Ui0x5Bkdc+ZLKBr
LyD9I3RR7OnIi2rtgozvHdaa7Fz2DmoNDVn2rzJaNIvaJtGcW8KwonQdZn5bW/Dm
/ihoWIAXUHrSlwOzOTK6uDEQtviUlRxVVP3uxfNNlFU6scxtoZZbInqY5oxDGpRi
jU7JtSTJa5jA/L5IdZFLPq8zOLY0tIojZ6Wfo9MZAz/Y09B7NUORcauqzyKkTa+7
FV2w8fUIETCwCb7eC4S2aczKdhwIRstLFoWsv/5Rv/gUZwA2e+crboFewilR5Lw4
OkAGqjHNE5IA2135z0hKlwRsVJ16A4p5CWUGK6RMnwJ0jNYzwXUf+Rmhrxa1Km+r
StlbiZ2c5E3XK6TQo7jkRfOqTeWBFMFI8KdE0X7Gw4OgZzl4Gi+kVrHDgslKRmpI
ieLncxZzp7+gMWHmrF6stXyZGLv1qH8nuBP67FoKo/kW74B2+jCkyIhpyfsM3eIc
rImjb8Jbst/zebhLAaBERgStXPdlG7iAXLqKXMgvb3QD1+gV427A3TxLf7Gumk/y
Q+d7zWhGeTn4jQfuEZxU5zSZbGOs10wUvhIRGJR10JBeRfcaQidZS2AGbZOoGWH1
rG792HkijopM+Zk3pZpA9sxhANT6OchGiglOp/YlGJgo0lWUuBdKgZfFz3UQfEiw
xtKrUGZ4K9FsWI1nZimv4MZciq0Bx3Sx7bEN1r3j1kbrEo1C1CNvlaWixjgV9IgL
Lf8X7IsrVD+Bcwa5Eubshv1puLDvjR17hz+kl7tSb5oLplQCeew+waELzVEMhFdK
/Y9a3inSNJ3p+026oP8aVwNlz/HRHLFQ7GIPpdzeCHTjKObspjg5ijp+Lk08QG0b
zecMAj3z5gKV91vCnwwXFxl9PpIkTp6CZ/ihTsR78pv+MRblcWjheROtUae2q02F
fhcH9G1kwPBFI36rPpPjmPrL+7AyjK1IHnA2K6jGvbYqrhA08EO0iSnzvgN6QwL0
NANvQ9lE5L0k3atVyNhtDHhUQywFG3hp3uFGdxv0Vn0R8q+e5kSZDzTOvfzlfLh8
hCxUdIU1juhDL4n8Ne9Xik4bPKU/IctsPWkSCWcyTqCsyMQ/qeqZ0IRZlyr/bpXS
tcev7DgB63189OluBCWst0cHc2i0LmqUo4FGQlXPd1OgretFwA4zBfrRKSlBMSon
qGPBCZcXmI0Dr+j4yvxDeXDMmTflSSqdISxuBHqkf1k17VA5JcnuxjkaNHO3zJff
THF7iZmvWAWDeMOeQk54vmK9B421kkTox1wnun9Vavr24Gz68s9th7J1qHKUqVtQ
kQoVwjb+SgmdTpYSbQEVke4uS8TBShAKufGmZEsZ3rWzi5plDNhK+1ElMEh+kQrV
H7SDWrNcWsioRkRmHT3PQA==
--pragma protect end_data_block
--pragma protect digest_block
Nzf/asSG0t8+RveMYuxa8dNp9Uw=
--pragma protect end_digest_block
--pragma protect end_protected
