// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H-?G !$C<FFYC L^XEF#4ZG0;Y9'.!^'GTT04UM9$5[FSP^'H[Z(68   
H,PU3TYU<GLW:%8+#F1WL>8,D%KD;<9;GVW)= JPP1JZ>A8UF8"V^#@  
HV/SEX2U,+#G,*OZ?Y(5Y3-ZF9VL/"NY%"+Z.N1!AWN6<= G@V;^;I@  
H2#I5Q;L8L9J(ZHH=Z6P4I=ME]6+25$_HC3D?D:ZNXWMJ7!$BKP5ON@  
HZOUQSW JVA;N[:V[I\5Q^J-T;+T/6;NHJZK*4E!Z"SGS94:3Q!--,@  
`pragma protect encoding=(enctype="uuencode",bytes=20688       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@BG@J'!+U#<3-KH/Y-,UTXK0[$@N+Q62.B"8H"&\?J,@ 
@@L)NY;%C\\Z_CM_1#8FFNZ#C<5)=NMDP1Y7H!@L>#U  
@ 7"7_1?%%U6O=M5J^CHN$0=<'L/9C<]'EPCG$LDWB?T 
@?MCF$W]JR[D7+L"GG',>K-JN&1+\[4]UZU3VP.;<?BL 
@)L%$^MP(38WG=-T\^ER:T8!IHR&)]7U9-Z%8.T@YSXL 
@&$WZ@,@"F&<(D*Z<>!*B4Q/H2E#RK8'V?J!0!">AJAT 
@1"*"[1NEX/<'URLNFDQ.Q#1?/[O:VO(M^FZB-%U(PHL 
@'\DX/@%3O]E 8T;D.;5-2N>SRM>1&2Y3 6GZNK/>09@ 
@/^-TQMR'NS5FMC,T8)KF@X/=/U>'7RG U5>SEE6(GR@ 
@DU0, BP;?I8@*M:$<'$11GNUMU7[H'-GQ,[L-J6\UN  
@%23K1!D5YQ,&$]0D-";^D]F9&K)+(AXU8\!YV%^I*;H 
@;LT>/^.TK@B#\0:@76,(L^!C-<A.!VY_<M\A!U#SW7T 
@/_P3 +$,L]WNP*6&']DL#!*.;F)%V+_TA_/MFKFW@[< 
@VP"(Q>BUKC;OJ%VI"1S^4 5:G@&-\YB:T0D_\;QR&(0 
@6S@XD"T:57O<*QK53T@A"^9!:#;(YC79+WL3*50@J 8 
@6R<:WWM4@=!W.(PGU$([1OM\[5-F^<P\ZS7:35!U13X 
@)]X?.0 391 :L!/D4DC/)*M&)I#1S*U(9M("\KTU*,, 
@\?0"HFQXQVZ)@[[(!L9&CF%55EJ/Q) 2(@XA[;AJVB, 
@J4 3F @ K*XD-0-XJ4MG7:I"+T[[)M1'5V,?0<.7!6  
@GS;("08(9D _.(I?5I**"ZJLA@QTZ2O])DCQ"A( 9H( 
@U*'GW+#W,/,S:&4&M[74#D.3ZSUEO?JI/M>!8(QY[6( 
@E(C.+D2<]%'2XFX>U"$8&P]>9E$8T_P0ZS\/\0^@82P 
@=>B\.8YR)+N7YW \Y0RWJOS8',R)L-T<0<XP^3_UGM8 
@$FRS(,*RMT0^ H54\;B&O:SLCJ9;OPQI 8=R@2X1[_X 
@&_MR-IZ&7XY%\$;?OYQ>$FX"._!?R=+QWOU@&\2'B^H 
@RRE<"=_DOB8ETBC-'( J%H9_<)MF@L+G+Z8(EX9S\NP 
@(B&L8=2^VN@)QR ,[8Y'[*FWQB_,>-X"+S6:;M6T B8 
@?050$XC,3K4WJ1S+(Q)/@@'Z11+%8H[EK2HF!/)V1[X 
@FZ%@S?YH"G\Z@$/8Y =(5-.AXW2O8CKG]0NN*;6HY)L 
@*+1,PP=H#BH<(MGN0)^$AB>-4,A&1OIM?>@_RMYU'J8 
@128G@$-[-@:0;FK]%%A7]$VHKY"*HP/@GC+2/N$[MK$ 
@Q^W&@"47N A./L?F*@!4BS];+P$.S=R5?JZ8,)$6PBX 
@11DVX02:3B5]MB#P.>=AFN##Y&3.REO$\2\1&J&=[O0 
@2^.)<,R>6G- R)V,]0C<I4(O!QR&_>[0MA4#'2"[LSD 
@JF@0LY*=NN83[>A02(.Q:;N57#KY\.%AF62I+WO$(5\ 
@AA,<8G(G*@OY8*U5ZX!3I6UE!=_MI( .<-5G^(D":L$ 
@J?>RUKVP/7!+U&MBLQ>:#87?A<C/&06K89<^V$G84/0 
@Y&QA(,6#DG5(I59(#2:(EG_)YT;"E.F0"&W+! 'A^^@ 
@M#*OG78T"+K++BQP1SAVB15OP4JV=K:O)IE1V2"PP\( 
@"1$W:KF=$/B#@L(AD^(NA::QNU(6KN7H6$%EX#]AE@< 
@^NB1G"2ZHX;F>MSD:>[NR<"-2YF) _X$E/0ZLU*B%BP 
@<X\I;Y]GPC1Z3]CY E875/]0J9%('^4+3:\Z1MY=X%P 
@>Z"GSTB34E>=R5R7@54J76F3X1DI><GU"=!!<V2M =P 
@DW ;P/F.>QO11(%_/(T8[H0N<&'!FR!,\851^&IOQ6@ 
@SP&Z9RD<HH&FBR@<KC( ^5*J)JBX#(&>S[M8N7R!**$ 
@%87M@*"\?I,Y\"\89!NG0@>:SYFC?M)*Z0GRMEP?ZC$ 
@BD#K[[D46]D*9_XV.#J7XHI&PUEK(3*VBCVEO%!.A)\ 
@+71_MYMISX_WCSWRM ^_@II/7&B+W2G7E5FW0,N1*XX 
@D_O!='VX;Q!UQ64"0YCQQ/G-X5:XM(U/Z_$1E*FDJ"H 
@>/FAP1J6*D>/PC\2O-ANV"71D=]E6.3\^C [N*>09;X 
@,FBZA'4N[Y=:&=@XF\D'I*=\3T$TQ',0PFC43)T191  
@+S,K 8EW[A@VJ<QC ,*T8ZCCS#,%/"82CZQD,1B#Z!X 
@\S)Y7B4#41W3!N59^W61,M0\AL&<BQBBW_L748_CJ@4 
@1+IJC;)O(W/6]'5KO2]AY7G8QG]#DQ3ES<KFC8 N$]0 
@&@I-M!L[8TR.@YU*15\H=27O"C/0AM\B'?ZOJ)(A^8( 
@F27\W3'^'(TR;/[LE,K7]8PI\]M!_\O*S-UYD>?K@., 
@_UY[(%]&X*C?-V/$T_OKR'L'P_6B$9B(<H#/%SF=6@T 
@U8QFFU>G[.)*#OLFJ>[7S9>.Q!2>X(N43?\$.POD>Y, 
@Z=R+?<1%K8XUYP34/;M(81"6<0#/.YG$;>_-6Q]V9:D 
@M%[9CEL8O^32X-(.[I[A"^6I] Y:5M*ERJ?=7>X$7JH 
@P@2\UCZ(!>W5T9U5?0@_5D5<_/KJS_FW.HBSL@^]+ ( 
@G+LJ/NU3S*YIJ=FV76(Z )# #'3EV9-:>OY/MH?T6'D 
@T<(>*2(6-^E&Q2$2 4RB:Q10I[J[C8&79&1DQ,!4Y'@ 
@RK[7TS3T3,:P$A\,K&PQ]1/OV&>_I\PZB\XVW->89X( 
@TGU@),,RIR9DEF%R'7P!:>J#O57"-W'>[%(0"F42!JH 
@($#$BC,\XXYR+5'L U/HD,X!1>T2?P8K>;)^^>=L0"H 
@5$$6%17&')(N0[\91I,HU:3&WCF_3RGC6'.&NZ9^\O, 
@\;P*.4Y6=>;_%9?6CE_?" F357GG.E%5*I#-V7<HCY@ 
@.Z(\LI&VL!Z;2+1Y#,<2"D#,F^R"BPG-FH"!L-#OC", 
@YOGCR0,@4@;M<%TYE6?,+7L,T.G82!+2B98PXKO,YN\ 
@D23XV0\WV83V=72[CE_)EELQ#'-:>GRN]7 +#2\@/+0 
@OA!W4R.9\MN4#NP86P:- 8AY*OZQDM+'>N^2'QC),/0 
@MML58OS2<EKMF9-4IT['Z<JF9#+YNBY.$AGII$FTFWL 
@H3R75%E4#)'WDS&JK?^I>&CN.2+Z?GD+%ORJ7_V\]S( 
@5:A>MG"3A.,'$BQUW]6]$58*#S;&-CE!R"G1L^BF+DX 
@!)V:A_TF\0[%E$C3;*>6^Y'3[M":T[H+*]<I\+HM)IT 
@I=5Y;Q]^\2LF:P<1#QS+--+?UR6$7F9S[M!^\&;SE/( 
@*':M;YPTV.H',^M"F1]D\!MPJ%/+_EK+G):H2F(;7U4 
@+XCQ^UATQLS+3G61]5VVIZ?@3CF$[W(&PY&]-M.LJHD 
@86?FHOA&4HTGT)9T?QB';&/67>U"=7OU!(XI*+?X>FX 
@:-,&/<K:Y=O,5&^)R1QK)#L@D,]HH$N'<WRO8=AA-C@ 
@WGFS!K\YR%0@&X5EAT?AV1C)G,HM[Q%8)R55>SOSZ;8 
@DJIV3_M>5H+Z.0E7":6ZDS4PXR11#"F['6JQ5(B#MWX 
@Y5]M5*$87M38'9IN1F&DI@RY/J:N2=4L$$=<*C0(*A$ 
@^%HJ?"*28S*EU*.Y3)H*HC+&D07F(*9&T6(T)H&E9X0 
@DO1L#ZEG(F*$0O0$",APSH!@D)+,D$<6=H>6U3J.X50 
@MV:5\%@7%5F<]Y>@(A\*YMV%N\B7D8!*K/?D57YX"$8 
@HM5>N&TI5VP!B7G<H$/,&LA(,-;H()WN9EO*MKR\F\P 
@6!!8< PAT@!$:^C6[8^,+;7=\KFLM@2V$;2G[PMOMZX 
@A\3@4R=9P 5%&S)6R)[\4^Z-;YN4.]NL^1%05YF/X7  
@4'F]9-L3&ER^#%0G<V[G! ;L'HUVG8#"8FK7D*IA<C8 
@X5:9":8\(7=Q3O^1I:A=:Y0^*TAKNVBEY>%43]6^QA@ 
@M(2-FJ.VD$02+B7+6&UV^)1Z^K'3-54,TF4RV8*W82D 
@WVF(7$FW%PI*><OQ]]7 O8\!A\JN&DGC<!EZRJ02G$D 
@TFB7 GJ.OX_.JW^V>;KUU>2"4Y5-%R0SJQ691E&DNG  
@XPXIZKK>M1B/;F.Z?&JB@,+I\S@5&FAF9-< $5[.QB( 
@\1-E(2N2;<A:D2'I(TC]3[VIU.LP[6^\9'H_#9RH'&\ 
@X97NO9>IWK'IKOA"4V)E4/1)C$%)6420XM.W;_9/6)@ 
@G4H1W71JC%<NR2%/8HFC"^R>OQ8>3_P[/9*NU,'%Y^D 
@,HC8WQ/[+U!^=-@B^*P/;IHYF*DO<><C+8Y82"<IEJD 
@0A9GE=6(@CSQB$LOJ7G8?)879D46D1MX&K(8A:1:JO  
@J'\>(F_V$,0A_G]/O?-D;[Y6RLKS%<L+BWXX:C97[4, 
@.(W7=\)3)=RY.U0+\X*J@>TAD;D!\[X2#A49T)*F!6< 
@T<4V?Z."AH$I;27#KR,4X1^!#::GD757J[0+$6G(Z:8 
@J=-XAK-[CBO3P[/S0HD\PT@*,I1SM2]\,;7V#&/>#"$ 
@AW18MNZ9$'+#-M(.<'+!P&JX=!M"F$2LH!8A)L,C2Z8 
@IJA2=K6H)C@9J;82%7Y_+H5;,,:K-;N83N<\O([ND,X 
@7<,3/E4H@\C:E$$K%SK)/Y+E'N,/JG-4<&5S/$]U&I, 
@R2 ='Z%O)2ULV^U7OK:1_7+]A!=N4O<>5AT.AUQ63&4 
@-7I%_.XV%>LVQK2#MB-L\AN&<-PKOC=G622/+RG,/L0 
@E#T:B/8W>7'P 2,$"2T">C6,T7^\!2\KP[W8)9L4@]\ 
@$&MI1SOD18HKTR_V";): V!H3:FU$@213%TL<!+#\10 
@YMH)MD&[ZQ[CK'ZP2:A5[X8=JD$S.IFI<7,D-(&;7?$ 
@AWO?7.\F@]X2</22S[TM5$1>LDR@+(I(DR7_O_T1IET 
@1W[D:301:H]O/7L;]LA\YS #7BBH%9B'N-KH2Q2:N%8 
@G77[DK*F\.P^G?HM&$?PXL@J WJG6^0 T7?E>FPS1GX 
@,!,_;LN.MK;.N8H %7<K)#]B)9U82+/?_9D(-7X@\7< 
@>MT]$^\&HCT?(IR1RVP\+M+XUH-U4?BEK#<,J_]C8:\ 
@Z"2>X@MN[O4R;YY,@-UYC>80%XSZ#<AS?&-5'<Q1)<4 
@U4=471R[P$(J8W3]-GOQS#&)_WO8O0I4> *$[T[>C&8 
@L/?B&ODT7;1@U(17W_(C<^$"1+'Q(AA;=:B'HZ0TF*< 
@*S,WHL4],OP2'2;Y[FZP&L.F*0)VW;95-.!3F/+=3\@ 
@^A$Y>FA0B)/O&^IRB1SC4T(8D-:71P;H\V%:2_[3]3H 
@%6Q_:/P$@STE[\[73:"2?>3JO5"ANP%#*+ %>KMR3.\ 
@160$#RCK?BGM!P@M5]KELEJ,V8,:RH-D+"W^ZW_XV;  
@'U-R*'8=5>@& <4^[QB;/.B;^1YC&J*%6F 3:_+0?/\ 
@RE-T (@,ABB^F!%A*)'NI+J/T2(3/;NRP95*+R6H<U$ 
@']T/V\\*[2W>,5\066:X:(=24P?0 'N[3$9C\;-TAEL 
@\.XQT(K%>(#]:K50P2Q>Q>KR]9-L0,KH+)TT>F!LN$( 
@,0O@T1*=%M5.4IGZ"W"R/.5?,[J-#_]E\E@K=T'P-], 
@H848B+K/B[Y<N*C,PAD@*9>)@+![VB?(HF<4PD5VT[$ 
@"T62J,Q/3>OWMZ:4,?OY+>6-N\0BB;T-_RE!"9Z+78< 
@C^^2/9R<V<F0ZC[VMN('0GB$*F#/+95#SQ[U9^#'2"( 
@'0<KR.+4O^>:I 9;9Z=?.<!*I,O:+'^2.]0&39)H3>0 
@P?;P/O(N]*+SP=ONZ-:X4";,WFYWX[A&]3^DQ)##(3( 
@&;)#'C8,T^:=M6KPJ%)7?2YL9T<E&J#'^!?D'C''\6T 
@(D#Y,,?<1IEF='%2M$MNZ"VHBE^^M$G4^DSVP!&R"!8 
@QHBR9=28N9HU$UTG#UQFT^8I@2"_"^UN=V81!58%-3( 
@Y^WYU^>J\?G-LT&7H\KIWIJ2?J&C%9:D,4X,U*+YYG4 
@P\(PH_60X.?\02;>8^%DIF31X<-GKEK]TD]95A6CWJT 
@LPKOQ.^*/(;F@V_'DI*;D+.,7SW[QO =C6$=$WP<PY  
@T653]OZ8*Z]=2(:AV8RRO2^+F0-V5D$TY1"> =ZQV@@ 
@<]30T*LV(V:^1+$1@9*H+1&FV5X)/F;-R$%.BX%_CR( 
@40P\#I]G>!.F&4$GA>KJ6Q$:Y!H@@4&)\J\G6EG1(;X 
@*?:9/6FKT9&3OT/TM^&42!I-H73G3I976D99J(63?5H 
@(3'UD$IB?3K1VB^3K&#N6/73Q82UW:A8K>XYIJB\Q0< 
@>87-!?V[*+Q&UJKXJN-?65UU>0%_^C]X)SEDK4ZK RD 
@>T0 =TN<2Q;N6[*E0(FO]O(5?2"C-*B0%$]BI:L5Y]8 
@REP:W1&IA]E*0LU#JN\/'S-BM$IM^^'%$CJRLL$F#XL 
@)A@7A=.LE;ZIAB.8WVF&@]Y2^3E4(G!MG>! \M3<V/D 
@'2S<]R,R8"Q2&<[DR$PZ(Z6VG(=P5G=',V;^;&4HW<T 
@@Y=QUBL/WI+D<>_3<47]?S[3D=NAZXTH_, AY"" =3\ 
@U+/EBC5')+&(OVT/RR75&AK%;+7UFQ^:C_0H.04STLX 
@&E"B_9B9]M?4,N _/QQ['U0TLPH1F-CVP9AM29#2/>X 
@=>*4O6WVXKRG$664 7L5>74KIB)\4O>L3IV^ N$W(AX 
@ET7-P,\5KR%@Z[MPSZ7'*KB -S$P=SJPL>]QFY</V?@ 
@%2#];;F;->4G?FPZGV;>'9/DQ_\TV3M!1N2V4@2@B$H 
@2.:[<X$J+$%=M7&PL\84&E <K\S !>HS\]3X^^5QPJ8 
@>02]!4'PJ:=JCZ[6\[I9%#E%P7?_O/6;VYX/AK8)G$  
@HZ'J 19'.9]'\F$AG!EM"9ZILY VD+%MPV?#V#G*#5P 
@H?[>O> T-H;EP%,C3]LO"K@#7/R[?WXV@R2L/J]$*A4 
@Y#W%]8NK01B8^;)GP7V[=@?')<%^7+]!(ZT]AJ?\_@T 
@"W"]CP>]R%!-_<)I*4GEV0>8ID8P3YCF!V\.;T'Y;F$ 
@3S\,898*(VGC>W7[I[, &A)(Q,9L[AY<>]X=3)\C$&0 
@O%$F@JBE0@FK@-@>*C,Z%*PJK^C25A2#NM>3BXIEB5< 
@/=*60 OY^;@0Z54*BNWJD2@5I&_\YBE<GH3ZOQBPV*H 
@_3=%F$*A]+(SP]RSK4 WH\,10/8F(<:CGZDK;_Q:<Q4 
@F:E)E_A;IP"7?H=WT;SGR7"+@Z]#F]!AV)D"OE%.^?X 
@)I90XW4'^GP68=U9% O9AO$?/*9E#RL(TWPM?9.*6T< 
@#23:(["R$+2V[Z_GA+&9)D4S!S8 Z@$A?UVP02E[&W$ 
@<"M,LPCIL/06%)(*"2.LZO1M#H"F ,(LWZV859]H0&4 
@NTW-]^XW+7,$972.73XX>/LIN=1*&\>'>ST.?PA>UN( 
@E:,KZ.M41BC:!71)50YR'D&^H115J;P*[E1I3Y?4'=\ 
@DWX$_JMMOF?,.$E(;JY#3312)Q&Q^T5];0R,G=VZB=< 
@\.=&:SAZ.+<BO-3PAX>M(!8W,NA?RY#M-BP(TI:DT.4 
@870 RSTB%%L[-1W;! P0Q=KV %J;:S%B=*ONV3+I:<D 
@93B$<&:P$=TDPG9R+X#:19QN<F$@J^XX]U(/]H%@W]@ 
@B%%;;=CA('\4Z':X;@I3)_+!K WR*'43HH.)R 15Q28 
@>9O[9U_(=:P=B $$#O"2B.]IAO9 ,T\A)JG^5MB&S3H 
@5!.EN! )7%WXRG_>^)^CQAIO,_Z*7E>%_=-0P.7":<< 
@5^\]$OH25M0JR8S0/<SWI&':Z[5( H*BH;J7D);X_5H 
@NI?'=#_Z-8TI73B#J@-36?>3$INH/0F+!"2QK<P?E]D 
@+[XQ$Y[(58J!&)<Z%E[VO)$JFV2=I["OM?#Z%B-WX=@ 
@02\B44[,LZ[=_RKQ%\UGHKX&,5)GXSYQM4)!/S_K&/\ 
@;QD66L!C&&D"54?Z#F%R8<& /)IN&!U84WGU#E?K9WT 
@V^]M6E%S;#&^-!AD&Z(HY*0:9YUO]%]&_6--,9T<HD< 
@+3ZYPC:?)U%G&<RQ0=+(."3VS</$!*N7/A\:H=GR[_0 
@EZIVS XH,9N$)FB,=NH<P0O6QA_AVE90V+!%<(E(K@0 
@)W]S10<4[-]N;[WP%PGX].C0+YI6R5R1V3:S7,T*SW\ 
@(EJO"WB SSO<DQX$,M&)MX&DP5,HG-UKD66+L"Z3G-( 
@LT2670AOPDZ")=O"<Q7>D,-K7UDA]_XB\UW?(-2AMIL 
@4K1V/-=]#UMJ9"F6KOHC5\+78R'(5$$@L-Q704_ \+\ 
@*FNUK?XH,F1R3>T/^V@*/* \_[S(EO4T+KO9,]4V-^L 
@)-1]V;R:T0>1A%6:GL=)W79U*1Q+-;U1K$]*B++@UO0 
@?'RWEFT 3] BL,D(5((3?(Y4M5%Z^B4) #Z5B!#&_@L 
@$F8$R:KQY)R1./<";2F2EJX!Y]"YPQ0 R7;)XB+'_^T 
@NY@;VO-6TE\BME-T(+\&N6$"W'NI>-4T5'UG3N(::HX 
@^E( 0J6'W&DG4?-$5Z^P9WK0RIEZ"4V?>F5@5LA/SN( 
@S<&*H(B^>[>@#["X _<SM.&$D-[I\9_"XASIU*):5+P 
@RK9R&2X1&"'K)F<???=YA 0[F,+ ]=?&/A1,>$$:#K$ 
@\.6K\EZ?.9% R.3W?9;W7V;*9DFX6<7HJO6CIM)5(@$ 
@[5:L74!_DKZ1<R6V*85R*5OH'C:)"9M$F.N],*BG63L 
@U>C"FZ?^8O?'O3]:_-TG29S_.''!\%(T:Q4ZLPW)P)  
@KZVJ,(?@QW5%IN3<W97Y8.,?M+@@6#+=@'6\9K+#AAL 
@TU7V,=+LJH:4HPO*C".HPFO9'%504'SML"4OTI ':PX 
@9";*3)@0W->:R"\U,^)2/[L ?"EI@F3#04_GT$@> QD 
@$_::UJ$@4\NL3+E=4+-"CA1#?+7C"+XSR.MTFQZ0HD< 
@0EU^6'<4Q$-V+IR(#]16?1RIZ7OB]U.,/V"-\4 ,'*D 
@(&_N=H2S29^SZ&.N+U%AWSY6M6NL93+ +W.5.4Q-5JP 
@M<<1L97:0<"?9:5>2"#2KB018\K(:Z,7:8'6#X4(**, 
@2'[ ;:#A3_N>[3\_\DWBO^63:%(>GN=RPK5[P;W44K4 
@+V6N1DV;T#RQC>&?82'#!69^!4ED ]=?.2[@Y:L)T68 
@D@E! 4YAM-CT?PEI,FZV_D%G>/9[K6 =EP<;B>)QQ2, 
@R1B9/3F=ZQV/(1>\_H3(8J4O*"=2]AJ1Y=_XK=2N!^8 
@XSOSP]ZO:Z):O 'OQ#&7%+:V(F-/:BY5(% 4@3T70   
@T;^(F794TIPB>5MXYU3;R913$#EGAPO5ZZ9E2<8':T@ 
@+I^"TV7##UHMP1*N_^SCWLIPG\NR,N\KC(G=_ZPH\,T 
@+$T[1@?84F/?]?93M7]-4^WCH;J"R* LB4JE=,#\:^@ 
@O(H,@9NE"?"*$G4CZF[KL>OH':Q..*5!Y,(9VL8MF9T 
@DS%L<XVCG3RT\[E9Q<>60T3@%U[Z]HJ=]-,IM=T'$&D 
@\2KLE#4D S_OO]B?^Z8A'</3[A1;H-DZ7GJF%'DQCF  
@QZ-,HPX'+^;VGANZ#!.EZ@D-'MW]ZGI81_A.Q61,&X  
@/5X&B/$K:MU4L] 2 HG![$8$'\).P3STZMC>(:.R*)  
@T?3E\Z%DX6T0"*L#?>HU'QI=K( =8(A@]X='.NS-)W< 
@^G KS_.'%%(FN)^8P$DF-ZCWJD=$$70:=DK15@.LVT, 
@&!02NXF9V@?)94V/S_H-&X>%Q!\^N5#1 ".H<S9N?1$ 
@EZFMM[V;2>B(0U**9H74P0-2HDM\7IF5B]O2F$C<+S( 
@^STIMJ*/W-X4ASB+;R)T(SB/9XX#CR,&UM8CPC<CAE4 
@>ZTM^?'*(%AL5-%=0(R8@2.'6Y2%=*WDTSJWB!&93WH 
@9I!FAXM>T+/YEZ<=U3.C>!7&)X?C/9>_?[&<2+%CL@4 
@JEN_H]F".L@7\Z(42FF(AJ-GM?'#G?T,G8XBDBGTY-0 
@7!F'"AX/[:;_H0' 9]RL&BI9CAR6Z[8H@LDQ9;>/="< 
@J9W+CHIXX+1OF(ILW=_C_.$A:O@V_WI<E;HRE3V3D6$ 
@;'(O)EM TJ.#WOL[Q>X1\7\S9;&4K 02_Z[6">,7DZ0 
@%$ P79#/0<3MY+:M&EY>,Q&R\U+?F@4CUL SI5 U>(4 
@WJ1__/HVC8M@3!,FIV&Q"WY@C)O'^'B<?I^7_N/(UJ@ 
@;?F+D-L@]:F(Q9"E$!'DQ>.K1JS/A=E;I>.D/N8.A9L 
@(KLI^W^W'=XR2<$%08OR)=<%C]/98$53AVTN,[07>#P 
@:Y-R#_YC_?.6YR[=FH6[]@"BI KKU:^NQ*QGES#Z]4< 
@]HYZLC(<A\?8$5GX)VSUF($+;LIS $<"H<_:^?HOEI$ 
@S2W(/SLJT_Q<EW-:CW7D)FV[BL@::NV&VC2\)]W[398 
@!CXG="E>^56A[/V^@5/@6YC+S;/WQM@*]PU*@?6R.0\ 
@!X*[.YHTX\,ORRM'\BGKMR& 3!18CNGG<7FK]XB/A[  
@+=YJ090F_?&;+?V&!]"5A'63[T[%0\C!WY41,2O,Q_< 
@"<(N1@#^3%FLV(9&2T(:4P_:YSAT""27L=ROR>5HU7( 
@T55ITP:J<;%0F"92VU3KE&Y<93:YCX<::RB7FW>ID"@ 
@@#SN_]DW W'1-)+*_U\84_Z%]B;:H"*Q"X(9T6\')M\ 
@GHD9-80,S&$?U.OS!*W.,["*&YUAP []$%#[="G)JDD 
@*N*QXBU1(+%&'A@>A__-\;D^2%$+Y[&JH<F(LAZ/3$( 
@RUU_]UO:0_:+X>%2EZXW1R-XK\F>,5O0-YM%=*[( ^  
@0DFJM@A%XYKF)AH?OD*YURGC@..8LK\H(623RP9S%X4 
@\+>MW5YH0KA1EZ%Y"#<YCR@?E=-[<*K)3?S4039-IR$ 
@,_WLO+'G5%ZLH5:]9=W[$.AC=E\B0)Y2!M[;*7./DXL 
@RKP[S&-P8/Q]%K[DML COE3);MN4.@D*>[!RDZ8RI(( 
@TLWW+EEZ5M7\[RYY' 5^RVYSSG6%T5&CK4-N/'F?*_( 
@%J_4)R9?Z$$<[KR*;^7_&1ZLCD);EZ-KH[C>!G\](>8 
@XMBRA\/OYN&ZK;W^N<)U;!.^ML\6UNFG-=)CC<)> #X 
@1P@$2M8  )AT'R46C[+B4@/XUXCGA&.3#;D=)B4S&;4 
@$W,=7Y4(?465W1\UF#81)8>2=D4H'QG4SN6!CW(1:', 
@T. 6 +5W*)0 GD'=/U&@FM28/'K6Z270<C)P1]&U"XH 
@<"ZT'H :FX&GK ^&D\@7QN,>BHYUZ)Y,YY^NFSV3K=  
@57G-;-LP0HZP$:3Q;Z!R_+W)+87(02/L-Y=;D*A=GBD 
@ZG?89H\3#'YQ"*!F80BQMC5M%"P(/?N7^Q*"HNM^8TP 
@]/1L+M%:B5>*"]_Y_&>N3TVZ0<N'1KO5Q25!ZXL%JE  
@\CLM96(=J#R8Q:*RU*!.,Y(/#8PENE /[#Q\:PD; V  
@.1+5Z94DS&?@?G!LAZ$:+4U?O/7ODXE6^K4H/)XD8)D 
@N(1WI7RU9.RXHMDFE#9=%N:7&TMX9<0B>5%$X%I#<9H 
@G#YF?V!W,XFBQ)!+MIVZI[,TO9)NAU4MVD.])R=(![  
@P.P[;D(L4C1PG3:.3YN927@N V<@:X,D3R4:U<A=5&T 
@N:V,;I!MW9D^G6U.9,^!Q5?J;5=CB\=V61D/RM\A8OT 
@4H+A+G.(H=N@:/NQBW KH\C?).B;D.6FB)R\RBR^+A$ 
@R"XUX)H]SO ^WN!1/KNIW[.PSB=\,EP %._/+FWZQ&< 
@C?M^QPQRJ)KD3E0W^6%YKOBI-:$71$/U_1<S!OE7X!D 
@),$QV^2IWA6)XLO5S*9K8+^HLYK3.ZN8V8R$ S, ;4L 
@C)9O$8$W2I2UV/J<JLKBSP!)OK(8'')/9W04&/91\]4 
@XL&RY45;;_IP(9?))GXT!+0XH'-Y'BOH>:@MEA N45( 
@W?^64:I^-FOS?#UI#U^=(CLCUXB?VC>_IX:+^13.=', 
@&&2E!(H2?GO6 D@G+S<6;QBZ!O\LPP#-/)K8QQ>9 1, 
@A46\QIJ))]YWGJ%&>B3#6373M345^?E?)7 F'F8$>9@ 
@X5.Y]Y7JM18NDY9J/(HU7>(R8#R8#6<P28)BF^E.OJ( 
@P[Q)O;&[0EDUH<EX_)&;D$Y0T,#J P!Y)*WB<[C);(@ 
@:JN&)8)H<#G'/S2>'W.,\V=X<1C0/IE]*E)YE8N">(L 
@]O**QK+1^.SRGC\^SDR&Z9OO+Z"[$UEX&NSL-5'N]/H 
@-1(V@74%E(<2CO L.^OKAY0,FMT20-DE ^NMA][)I%$ 
@PHV/+D$>'GF3PME4(UFB#OCNP'OUG>5/L)Z6/>U4AG\ 
@SN5/P^5$UZM,J4=LJ+]5\,D;&"$BN:8K53I^MU33TXP 
@N*YR5=_;GT>F1N0OQF33Y#-#?7VO.#W"2':G09,ZZ?8 
@K 3_:A;2F%"W\V--971S(FM)K8K3+\B[L&!@>ZB]T@$ 
@R#*"TUY7^EY?/W0SL^5/FV)9?Q_<"++ K:>6;_4J!<0 
@TZ&C15($ALV('(]^ ![I88MHDZ=V###!A>/_^S]Y2WX 
@"=*Q4RKC624JS$N3D/A2VW6_7<%FUG3Y]WL(6UD48]< 
@&N%=?^%:WOTA=000\(HD0ALG.2$G>XX97Z+\PCS)0"8 
@ !AD^+)P/UMHKMD_182N,HF4\#2;W*[;& #*W3T0E6\ 
@6EX.Q:!ZLX4M =VW_*,087N(W 5C-18$+=BF'9L-1E\ 
@V$]B).XB>T 05A1*5!Z0'_@;U7CJ]#P-O*3.,8B&=$( 
@R"Q*7+:<N6W4,64(/+FQ_(AR[T1BZB7R?UY.#^?*[3P 
@R('J(U"#.00EIS:WYKE#\1(KU(*8V<F550<K'G',R!@ 
@E_VMNL;0<%X?.!O4V'^Y/_JFMI=Q+"'_^NMMSITCJB( 
@T:A;&.OS;?3NWS3\115!KJ$AI5S]#<9!N:>IGG&Z C( 
@ID_U_>-\Z<1-XDIS.4XG<'^C.(W("M#+X-BK/1.B/ , 
@("$KXW>Q!,V6NWVS1P8RRE^MG( <->#Z40Q[S:I$):8 
@OW4[$I/6'>E4@MS6AN8],O5Y^[&VBE(R96FI4)*A/<T 
@_+D?P17FYW0O7?V9(SZ);N^OMD82"/)*!MV62_]T_1X 
@\ER+VQTY_#0&J;2N?.M0+4LY\$Q-EMJ??\'MB5R-0X\ 
@"@+J*XA?,BBJ3OSQ0,OQN9"63,"-;/JKTCG4QN<I*5@ 
@*F^"GRJ-HG@7WDBGZ<@.C%TM/<1,]S0,*M<#Q@3<SKH 
@EP!&');X#>Q#%+R6&=\!M<B5$ZPLR)/PP:HIFA*,+)P 
@@V]9HJ"YM?)AL\!$M EJ*>N@D54ZX"Q\^K]FQ5S>9U( 
@<-'2@U.L91&=_FM2$_- 6WI--"!G@/(;$3N%F@\BVV< 
@]#H>.TGZXIWNFFEV(_J)@TD(YD%V1I>UL8KNP62,"V, 
@1?&A<3P(ZA55G$$W.&&_4;-[,-CTL'HV6WLVL<\TM&D 
@H$53:M1,O?-!VDDWDKV1Q?VOZ@?<70->7:>)W4X K"H 
@5>CAF;N:D09=XD.-KF+RDG!_X_DI#_4@:&PNL9OYR3( 
@_<U]/J6$Q=I:D1_H*K-3)8(R$-J_M7/\RDHWH(-%0]\ 
@J 8L^U4()N2F,=,5 JWY1'SNY-((CMH,$%7NY5%YS$T 
@Q(^O<:_=641[8U7T&@/FD>U#V#+UF_OD8ED,YF^1?W\ 
@KZJR6W?]92'#C;\IUKF\*H+I-8V9S<+\YQ-[0!Q6\RH 
@GG#"SPCLIO8;M.[JSO752D<9W'!PS0T]J,/8H^02C0@ 
@5@$I\67R!"HX$Y2'_"8'AD>?H)NT78W5SVR_3?<44[X 
@@Q;O\R#B5QA*A63W3:8_L RBHD,EQ0ZSY<C, MU\,4( 
@R]8+!.[POX0,3JW[3H@W4KGEYU-^K<3*XC&P*@WO"R< 
@]G-YK6%-CA@D9 [_$W3_ M\@*8U1B;))CVSQT=U));0 
@DZ>@T1NAW=@[6LJU='*PN- PGCWL'H/X*\!3GBP!?T  
@/"2)7,5#"^<1]:'CMHSL2X%!69Z;4;W,"5PO(]0GAG@ 
@M% &@5K[Z^LRO[):T"SET6J56S'\X^(+FF/=;\9(:8L 
@E_L.P0Y'9*8[_S]WD,&U#M")R3#/,"8[4AFQO;-;SX( 
@CB8Y/KF S.KN\26LO\(DNF^U$(/+U$F"C4I#IN[Q33P 
@;C\:U$FK1G,_[#U[, .ZWN>)$CC1WY@ :8NHF>R]G$D 
@P2$F%#E;:/.FFJ^(S]EYPI"M_05T4.0SI0%6D73.0M  
@]FR,S-I/6:UC)<:%M4*U1]C7=S,:C%I=>1A:K)**RJ  
@E+=#J1M4,UUKSG.#C=R;C+S(([6@L/-[0B.^>V"56/X 
@&)<L8AK(/%4O8\EY,@>ZNE YL'[M<@@F9X$!N$T!%$@ 
@7N^RW-C2T<ZR ?N_4+M[<II_%<F+:6!8OKZ8^BU+=-X 
@*WD$_3&.]3U*WPWA%1 J^A&X:LG:#ZO=[,U)K2,([B  
@WEGCN>".>Q3Q"4Q?Y;PJ49E?1.SG-UEH^,./WP,.HHX 
@-9C<[^\G78XGM_T?>@/("8+]*VI=-RQRWZ''2V!]2-( 
@I+\$A(!;=L-S5="B/%.-_(7F61FZMVM['TJ[DSZ8U*L 
@9;27ZLJSGH?=@<3+D[] @4X))\N^675J)'1X8()TJ&X 
@[:_CK[[^[M"P]&A7 -(I6JD*"MX"37Q;=7G--V)B>-D 
@39Z_!?<TIU&"I',7%7:Y"S' ,K$L? ]87\J@X0LZM(D 
@KR[+K5S920_QLV9LP5D()2L&5K&!R9IM!W)>?,)2:94 
@$->'9"*+-5L<@RY7F>YQS8'C&]OB;YA>&6B. M2CMT0 
@V.3S*#-<?:XAE#H&4O]1[K#\[R:HP@D.$[YNK%NOJY( 
@7W]=08K15Q+!OIJ-\/L89E*#$[=+9<4(-.5?A="ORSD 
@C8^*ZDGK@M(6-KJ!-9(\I[(Z>-@<P'^.RI@:IQZY@6H 
@SIA^ZXP/?JI;CWJYP$N[/,G<U%UPBCK\0=!\0TL/\58 
@/>N) 4 -'8_ZDR"DQ@XV@[WU1R>L%^RA5L>1O.\Q-W( 
@<#A\LDBJ9IJBX/ ^P7WDM<M46G/MUKG(=A%Y/&Z _KT 
@V\RYQ,X$5D&'?#%9(',N\<7?O4M#UM-F=IM@$Q %1&4 
@2'=Z (_]+Y;B0<RG;UG?@C$F]3#SQP_4IUE4'X6R>'D 
@T (P1!03H6A'\J*#B(]=$!R@DAG0G:; -'0K1!L]=AT 
@%\'ZVP LBA?P$(R($$'SV*< Q3"G*#JS&LJ1L'*ZGT, 
@) *H.(.-_OQ S8(R.! B$:K/8W+\)/^7T&F*<W[-^2< 
@O,.\GW"'F?M@R\8T5%)+$H84_%"Z#<._K:]V:#?_*OP 
@R+SKX.R8V18'G0>;;'KR;O%JKJ#Y_1)[]:\!D2$S,9, 
@'V$&.QHVBI<\D:VAHG8['X%KB>2C4+'("_4+VO^"6 ( 
@].DM5QH4\FH*P;P/?<$8VC.?R#XH/0S:2C;=]47$,OX 
@I!M>H:0XQ#Y@HE+5MG9*5NEB]Q>)+R2,DE-Z_,^$8,8 
@(-B@+9;\EY?8$VYX#.G+KG?J),"VFUOP.-G:8.(CF<T 
@Q#? 7@P-B)#0SP'5!C<RP]9&EUN'!UB(>N++(*_GB 8 
@?KD,8O,N>$X G?A1CG]OP5*>"U<DV-(#5G>GHB;?!-, 
@'6]510&G)Q:&I21<J6/ P;X(D3F*CFX9 \MK<!K=7X$ 
@PSA9R ***2D0%$CEIK,G!1]G?_7:E/XL]]U$TF #D+H 
@L(Y8!<>VJ[!!\UJB-Y3*N.'Z1-8NY9)344,S0W8KGMX 
@E*9P_[8;Z]3-:3JB?;*!,4,*";!-S_F80:>8_$]!+K< 
@=F(VGK3;$$=NT_!TRY&'78F6D"<)DW%O#! \_89RYW4 
@-#5<O](R*= AEB- ]120_VTEM!L2GYNDZ^TB^D\@G00 
@2P9:>?&I[AO"$(U:IAJ?FA_1X+%^;N;_.JRUI&AO(VH 
@AFS3]&)?)IHRPR6B/]G'9+]YBHD^B$9FR"])5+ 8\B8 
@[G'1$-Z\2>(3HIKC6LF;J7!IF\*!3FBP\_Q\^?"[_Z< 
@+Y&X7Z/*M+<R8%R^4'N0IQ7Q^CKZGB&<YU5*.FM'PEL 
@'!-5VV4B R2R:^TUV8\T*T>9L>*:6,?6@-8A)0K)H!8 
@"K72N_+ !F7N\E32XT3N4M:M%YJA.P-F6TXS->,^M5D 
@!D<AL\0#*!,(DTD]!X>1]?A#(E&/M ["@/W[.QRC&DP 
@NOU"06/!\L'!!P9C)VH\QUL&^9X.2B%2RT!4[WS,38@ 
@9,B7="@$+&?@+?>'B'N1U7Z^JXYRF_L&(%S+=A: '0@ 
@W-9AZQ9:7L//A#:UQ\7Y.:-G4T9BL!FS-D%0'-YLX.0 
@@WS)P42%%X)A,V$C+ RKFE0P)<TZ*_@@%-8%=@)X5?D 
@[*9>G"V0#Q!+_1(P$->T>I\+6%ZO7RL1UH@)N$W2))P 
@Y-&OL(^L@:.OJ*N@H5&JW<%J+'X+5#>S>-(<]?5HP-D 
@*3#-4NST!U@';*5S;-V08/HD#5)VRT;ER$(O[TKB7[T 
@S>1]I9^(KE#W<@#9^T=?%910("'V2RUV)0E/BY=Q-#T 
@9_-,4=>+?@0U VI-9L:B9&4>7K$+3 )R;K)K!23-\ED 
@B+I&'?9\I0"5PMU!*](*O# K^#&9H7/BW]#7E["SRRD 
@VB8C2S7TZH[:/_S U]U'KHF]357U+Q/F+Y3<NJO#&O@ 
@"E]ZT[X+^4BVMA9;8R::U]+HWABU7[K#*UL$?"]!W2L 
@SRQ8+BCR3!#Z&FCO M7WD4U7Z[G@F=B!\E$4(UJYVMX 
@JEG-$_%^/N?EZ-Z5#:T@YZ4T;B#E],]83"MN\QAENH4 
@F.[K6R<Z<DY<:X\6??&%#2&PJ4MWIA5QB?[Y$6:\'_\ 
@@(^L+HZAR9@@QZV\[?R^.&K,4%=E@,OCEV,0MO\S2I  
@J>-G9.#>07/Z*]O'U,*BR79%(0 W/HD1[81N"H0@_5D 
@A!'ACTIIDVKH*WCSG) OEUOO+37^$HM$JH"L.L7*E<X 
@VY(=^D'7'K(? <6#/,,1>"^B9H1XS;2G3)RO"$6MM*L 
@S\076!*NL&])R<K][-;'Y1H'<\W5NIV&ZE/"EAKD.$X 
@E8Q3*Y_J)27Z,$V'9HBHP\K?PK"&=5=VEZN0GCPD=7@ 
@A3F/KSD,BL3RA@C%X;3?7ES:+3\BR6;9,I8?R9KF' X 
@2\LF= (UK^9X;Y]C3OI9?,-8Z1DU)'$1BEHTER(0MEH 
@0_G&80X LVSY]9CQ1H>:%<^Q-\!S,_I\",:'+JR:HT  
@&_*8(QIYYL"*8K-J@I1S>LT0;EXA0K3BRSA7;"<QC%T 
@4IT;4^Y\7;@^*F0#501UP W@[H15;$I(VY>4MU41<D( 
@;A 3QDQ<SI33Y:>L8BIN! E'59CYZL:[/?!7GZ*N\08 
@;HZ?-Z:CB2NPOAVD8WC.L'U6XKXN]:N_6WWY:MC9/-D 
@LZ_+R*\Q'PXM9U>@,M@=93S5M#NZ;64$K&G?%;TCI8< 
@!-R(AAC0D6$T=X?V!67SK;"2)2Y*+#PJ'/.,[R.2WU, 
@%@>5>4.*V)I.,-+^3CC;KA!SZA@+HUK>F?-&'[;-0>4 
@FT"702<"9Q.&YK$'4K[D[H)0LC$P2 ]4WOO)[+JR&Z4 
@:;8\!^G\/+'9E5I2W<'<4,HFK\#61PP0>E^^ZQU?*F@ 
@YV5_IV$W6.0K69.P5#X0_O>R=:J0;0ZJZ*T4F /<9T< 
@<NH@FS<F21./XDUP#L! G3&Y=7DRJNZ\M6$,_^,G-/D 
@P7+?<]$S60&C8 R3@)A)H-=?=LG<-3B/%2?_<1RZ%QH 
@A+[XP,S*0<5[SR][50T]2X$E3R+^!3\<KQ2Y_IUOM68 
@;DWN=9G"D#_9.@S* ")=\8R747%LI/Q#^SD#.T(21LH 
@6S0BP[Y?\6IQV2K9 A"C]?%/@PH\ O^&E?N8TG247Z, 
@G-?JP'Q 4%X9<Z/8(XO6J.<&B8T=TH2)H0WL=H2-OGD 
@)'R3+,L=.M8,2F ZOO)7,RAYGW7(_XI4AI/"42G_K\  
@+7HF@LM-8L$4925:9&*WG_D!C/DHW#(NER*17@8GB!\ 
@&!+:G@S7:8:B!W4KB)FGK*O(H ?9B4U;1YH*A\TWQ:P 
@46[ZC2AJI?MX$V1O\ 0S:"257DXTLXNF@\2NLC;T/), 
@Z&*_R$<]=-I2?X+KN$DP 9\$1N,G9-,;!:V9K>*W-OP 
@=)8D%KI3JC,:4.Q9%>9JO\SZP7Z3U<JX8A7L<J^C3 0 
@XFE@%07_Q(XDUXV/U=)?<W4<WA[7Y::',&.2./Z@DZ  
@776'D$"*)^IPL7_$1?WN>XJ*[GIPTN7ZXV\9#]UY4!L 
@<0DG,?WC7OCXV=UBBN@W_2J=;P"S1&G&PF2#H;4+EJ\ 
@&? W*O1,67L,;5Z<U9*=ZV->( UED.L[J&Z?)W< -^D 
@Y(&C[1K4^]W/!J?[J[V(OH\GUA_R")E.BE.*8H'&6YD 
@:NA42P@X0IC\V@=3DVA-,*UPB.%>:LMGB .GQ.Q1GY@ 
@6'VJDC+^-O9.JP^(6_S:\K-15V1@\6/YP \%4:@9B(X 
@SV[^43)OPOA(<^9%TNL5X1!$(=_E]/(<C\3%*UZQX6< 
@WC89XD\B8<W33WT(8*B5T+? D 3(N01,B-W>;&^^3IH 
@*E?1>=(?_K$W+O>XVA4EK)!B_T9O?0?OK=^#^X[L=\\ 
@*^T["91;3-#[%:+_D*YF6,-H WF\K]%'HY+;-&A68OT 
@&.:&T6+;D $,^7WJ4NI(POU'^,#8:HA*WI$=W"XT1_T 
@=''9HZ"9"$H(#WJ?O2+W9T/"X@2A&UG)<7A0KH*;/:H 
@>H*<0W&'>ZKZ4E5*H>>_:J]=NW]N+5.;40+AP9@:]QP 
@=HS":O.U=G80JK+W,I+/Q#XQE%F&V^YDPHG-?+B5/D, 
@T)F&@LW+=%(FF14-1PDMATH_=5LBK/PRW*#?B]98@PH 
@2?]2)+) "%D(<<,TXR"U2V&[WT-1'?JGM1Z*^64NY&8 
@<6$&>^[N-5<W1S':M&5#R7%H-@Q#=WE0'-(I ]W/4/D 
@P5EJ9U#2W"3.ZKF1*@RCOV3[[FT6G5"*KS0Z!MPU!*8 
@&KT8(M[%NZL"+-&9.?5AI9IN;WDHYZ-&%EMR10R+[Q< 
@.78A71E)XA9<=-W1<5-Z[5$4*5U<9#%B%VO7II=4$7L 
@/"QZGI>'FB)?/GZ&+#54LB@3B"?*:"2'.=Y-*'0&HRT 
@T&N  'G4P'(-6*)JXC8,. <35]*V6I8Q6C0ZS+5MV:X 
@#I)V>Z=QCQ4$W9>5Z/^C\+PJKE[8/,";YK894N+6_58 
@8DE2G9$RR"'M/ (-"[_ ?/O)6K<OV)N@T]<#B-C'/-0 
@.EKSZJ\PS*/*J&W3<V.=?RX6_5/)Y3#1NU8VE&!D?QP 
@J'HKS^]E3;^W,_%5I)EGH(O[_G"#<G@^&^NFKHYY9:$ 
@VCGV@)U/KIY9P/XA/^<3#IK5.6SZS/<#"KF>*"WPO[T 
@6<'R%<DU33/3VZE$JJS:,(NY"#552KDXCLDC1IQ#V[  
@C=,+YSI@3K;%JV3R]=NST/EV R<FX A(F_98.V#?,Z8 
@@_]%1D3EN,%7;W=2D^,JSBG:+-C(8E?:THPYMCQ/VNP 
@V0\!]%GFAE5*\3?:BK<BKFS[R\'QEZ60:(UDPG/XV9P 
@T58=+PLWL=/_0EFH.8\PC(Y/&8UYQNT/>I[X]?7/H[L 
@W:MG@\E5F2V*7S#P2:'XS7,;$SL#DZ[%J1Z)O-DZ0F( 
@[,NNT!4'2#I /:Y*V0Y6<]>!CXI]BK,\W:6>'\<]N)D 
@0:#^2]C=QKJ&<^H.793JZ0'I$ZB[_OG JAE>.:_?ST( 
@R[?.T2CURR/7->LMLL[TXOT3%-*576?,'S8^4*4K[E( 
@F MTD(=1HE*LYPEH"WL'*"KKT"OF7W[1UOM?\N"EW*\ 
@MD"I;34K:"CTF(*<9A,@,,B7?'ZL$\+F0*?>!6>./OD 
@ Q<#N K_VJK2X:0.K2;&.&W)9S$I7%XL'KW@"=YS)LT 
@.13:(<0(%MHE/>;JV^@2DCOV5X_Q%)F8S5S#X(&:FU@ 
@)[NO#DF^&NJ 1+G:9@7.0?,\TX8UB2/ROW?T.-NV:A< 
@8GH,-2VM6*7W7MNF !KJ9D;\O%N>M!$GGF4(IX&468  
@9]ZANB"X\C"_=\M8U6SVQT3-A@8V[<ZE^PHN_%T-?QH 
@#/&RZ(<P^_1C;T%Q?8HML+= J^TQ ?N)=OX,'&N<S88 
@K7];<[W6;4,XWX_L(Q8IW!"FU^@G.S'.\@2)#Q[A3K4 
@&-7-/?9"=&&K340=K]-,8N+S&TR?]J>>2'SQI%T'T(, 
@'EDE-ABPMBA<-^L*N>NRHDI:S/?"D]^)R4+6:3I5;W8 
@YO\1IC%,O@0K\".$4]BS!^!=9V=*ZV HW]XR(\-\A2P 
@]\[D!DV'5CTJZ05!^+O'9^%#0K7/NQ@KFH^;X  >F:0 
@$"%GCE2<]%<7@$'TP\[6]0UK YN[+*I5K3W*<4SY0:H 
@G ($&H>6B*:/)"ON]6\$XKRY)>.@ME1KQ'OQ>!'O:A, 
@@!XH&'!$1V_U$TB#3%;@_"Q'9[G9OZWB\5TLKY<1K-4 
@X+Y=&32,I?&VBK@#H@?1+@Z7NC')*,JX2?EVXN=XX;  
@4+F-056 @B7.'[$?O2#\Y(.(NA>SKXV@Z%2X4=O5E\L 
@NK6-+R@U2]@'5F=]2)JJ^F-V'$77I;30E.0PZ;UN_&X 
@#O0."E0$O/UV5@D[05*I4*'6/O.+>@;2?#,.O0B!WY@ 
@[V24(5'@H5*V\^T )_[_P]%# QV.#LN\IR+0L1*]8+< 
@/=M1_2 B(&-^.:\'!U+)'_E>Y5/+U99;YZIG^*I*0&L 
@5B,-Q\(*E!U!:^&0AK?H[B0-U:HE^XD3* X?]CZS.Y@ 
@;[6EKGG;<)B5RXQ_K[JNNQL'8$8XI(B.-3K(]@W,%)P 
@>7SXT>R&A-0[&35SN?AF_";D3?*[3-"(=B)<3H![\)X 
@3X/%C@4!'ZD!/[ZQ'K?QM=_B7X-F?QO?P?6,XV<I>3$ 
@1 S6FR0?);MO&<5]Q!>>H702I&1!&16V* /K^*L KF0 
@)5Q;WN:OJB!DOX(I-F-V3). 4'X +S+]:\S7,[YSR<H 
@J-^@<?(.R"\IW?/;D*&$.RX!'% \"QK$WG *@5)3EUT 
@]D/!O*C+CP!5'@YG/F%%99VTN-K>!!1''Q8XC:@R?MP 
@'.!&VW_7#"4OYM1!G;NB^;:8KM#D&6"5ETM%%C$WQ0@ 
@73>9/71GT<74)\<C1)VU=X<65L^0WME;()MV=F'OG-X 
@,4=6,))5)SK[R\7WI<U=Q2)!?'ME>E]F"DC0>5GLPE\ 
@61+%= J*=';TNB^E#*H[XMK.;4.,1Y%8:*6Y<1=. VP 
@^H&"3KYU;7821(>H/4( K36@#LH0.U-\+>]4P?B[1'H 
@H^+8V4[^G,UG)B_*+&<2[R^CO %1#B#Q;N .O>;5\34 
@^-.N0P(>>7(9TNYB,G:PE-#DU--KY%)5ZC]?"YJ-<@( 
@2P41F(V5Y<E/5U3%VON8W_8]9RS8"BSNZ1V5TR:E"_\ 
@S377X.!DDFF?N:&FT;W]U.H.>TK[33E0ZD6YLSC^Z1$ 
@TP@2[;'*.9&^-W=CEP+/5<:&*9?E ,9"=-!*N3$8/KP 
@G6JH'O5!6@[6DI=*O*C&=]P=ZA%;CKQ42$_BP;FH8V  
@/-PVC)NC1"]]^!Q2&VA) 9N5\K:RO4MFN7)M7E=*>(D 
@:/F!A!:KO>@97#."3W0ONL2RAQQD\Y>2)TS<D!N"+Z\ 
@C['[KBT0'-(/\C6?L8XDXU7X25 +*.AJ5DT %3+5NYH 
@XV(D"G,LR_ M(+EFRO85U+-@AWN611%7+) Q\[HGOW0 
@U*"[=__YJ;9WEUX$,NM1DR^;QG*9%NY1]!WD5!^%(X0 
@VPT];:Q(R9^@27'KRR(P:SO@YV&MC^N$3-"Q_9/2-%P 
@>()<0MS,I$K$TLEN4WB*P0"*F?K/VI[UOB% _].+GC$ 
@KL('_E4W$-0VJ._3RW4\,;4Q(BZ7"@"[%ET(+$S!XCT 
@6=;GN;HXY#'("-6EDAS'GWBVW%T\Y?U.Y-6S7=*'TDX 
@8?*@$J&)/26)-6W27W/67+$T3#J/\1=Z2[#HWB"<(D( 
@<\ORQ(%V6C^J?&KG&0>K* W! EB%4"7SN&N4KR-3TBD 
@#P(N7',W.='=\J0<6,5<]2I@$4J[)XU0>Y&1)795Y)H 
@,ES]K*Z@!E1TW$FIR*9F?6^+ZQ@*"_6IRUS/'Y1PZ4@ 
@U%)<K7P?B%D0JP,A=JBD_*UJ9SI$\G<:+OE4:#;OKL0 
@L^?\ENZ+KI;Z/" >@Q4Q\L HN40DQ"1=)Y-.-/8Y*>$ 
@["(8E=]UK)=YA'G?1SH0"&D+P;Q5#7KL@.5(';DJ6V  
@3MK 8T/;%Z6/EC*C%Y=QM/6M$XE'*X8Q7^A"4H;>)#\ 
@:9464BA'RF-R_Q4\SSAN<C9-JC]3;]5(_8I+4H]-1#H 
@&FWGP%\)WZ"?:0*$ROE^/?$>\<L,D\HSCX5"-Q=$;<L 
@M,>E%OUV?H7^%-X+<4"H&+D=[AO-+G8[QM7.*DV+?)@ 
@PD6R3/>/'*'E>$#H=G+-ME?B[L\_6<4)XG/6G)#&1LX 
@G2*FK?O+;,A/9W'&[UFN?<&RU(@?X>ZT 36"+ =GZQ\ 
@H1]CW%GG]O_?%E#P4T?V]*TTZ\BBDMPG[[&J9N;O$,0 
@\:6RX133U:K(#5V8T$@TB[H?+"*Q[ #8#R[ZR:.7UJ< 
@A=$(]*G%-M?-+D_F;!+L0$].D?5Z=!$RL0;'M"!U4M0 
@!7+51W7OE0B^+.T;1ODCH\,U^C1> M.\*7-Y$,Y;9F0 
@#]&$'F!:7MM04N851-$@:X92K&VGIC^+/%D^[UYW+V0 
@2B*%T;*]BU\UYAP)I+:EAD%?(/>@5CJPJW#,?,E5PY( 
@4EV<_&VRPNC\RO5<C;+6#E@L^W0ONSN1E87@_)"I4KP 
@\I*W*"3J,6,5FF8KU7I-].K296:QTIQZ0Y\& UMYQ*@ 
@=*%Y"X\!36\7K<$CV'CN6$'.V]\&;+S57OG$OXA5:$\ 
@NT59:M=;Z&#0?)A'E6- %HB+]+YXB,9 ('],MX#W-P, 
@!) E)5<)P'HC7H"?]'9WIWQDG' =!\L- >&[0TZ1BE, 
@HO-I'-NZ+SF3Y\CY)9 Z?^RGHHJ#A>0QE!-T-$.8,_L 
@[YU>U=[XZ=<TKW(AXDZQ0U=>5H,(;:C_YXO^$+WF-<0 
@RY5R23IA]?J"3$LX^\#TT],!*T%LO:UDP_%XDO?0.L4 
@#AHQ<%>02Q;^>_9:13BXJ]1/GEU(&%)GM3P7-TSKEU( 
@_II/)]:BKNE8"6PQ[ZN0[H0R!K"" S\MWY(5G"A^Z[, 
@4,>WOJE7;@G,B?Q(98BZT%.*@M,0_8Z):VC_:A&^QS\ 
@W#\G E\UA'3(YA,)52(2N1W&-+D/1X$FWQRP:\M^0AD 
@PJ,.'Y=Q\NT*ANHG3&62)U0*<#[:J4<I^U[N^6#<Q$L 
@L9:F%40IGHVK]L)2@BKK#M/:6B1X.&-5G@*O%-C#O'< 
@[H6SW#U^#5,?VCI>3[S')DV5+\<HX69U&-36#+.T("4 
@)6K#X,D_2]X@O.?<FP'8X]& LL)ST&_$B\!#[J0!QE( 
@A?TO;6)M1[L0QUQ@.U@K$ 7_)I-EY.!!=6)1*Q@ CTP 
@TDG:92:2Z.ZO^32F@57;9$(EI[8VK G=-G"$8"LD;>H 
@,CC5H_\89CU/W,"&!]Y.W^0G@VIQB75&6</O0?;0Q_4 
@09-XU@UXO/UG6CVH^S%)O"ZO[^%87WK4'V5Z;<FU(V( 
@YPH)E:6 ZO&IL-9,';@[*OWIW!D)7%ER\A47>S&.;FP 
@O0F()Z@7J+)]^*1WE-1=[" 3/KB)"&33GV>J&#W^S#8 
@UI3&]G&6Z7B[L4(#37ISKH(+$)E@2B2>)TJ<X"1B2H8 
@\03=;7H-;&41%-]T32.J^U$O*0"7Y6!Z*>1T^B%1,:  
@S2.I\UZ<C.KD$K[DRLK)-^$:^!.855;0_4R\*ZK;Q9\ 
@.$";YS<\;X*7NK2&Y?WD8:+-L,O(R4[H'0)K);PRC7P 
@RKL>Q" C\WZ:B/DXOE:-#SY)VZ_DWIX:B7,MTDA)^C8 
@SFEY C9_A8P[P"$90LG3B=@+;(B!EFB$&[A8L-6BN8< 
@E>UWL&N0XZ&Q2I J;&'YNL_YGPAPD 7+UU<H"]I:"OD 
@$9?6VCOEPB!TSP S=;\[>7>.."T4_JLQT^RAKND"98L 
@RU_9]T4BU N>?PN6P=@,[IC?\CTY46H'ECG@IE;)4ML 
@HV/?0N17[[XA@E.Q>;$7XAQ-$5<[\Q2G171<V0"^294 
@0YQGGI0A&666!OJIR/$$G7T!VT6P>M* 6@\TJH&]?*X 
@*'ZO^&M;RXF%E4L3I?VE>K 8A#P)'5 4/B6\'M@MP78 
@\0,AVQ96#E9PL"'S%XFM*9;N&A=7'&GJ@9DU, R%-#D 
@U0(%5TQLPG_B/4]SJ&4;U!J4AC7RF!U;;?G7,9(IJ\4 
@^41SGQ8!AA*MSP LN6V-VIR_%S0<4,^P\Z!&E]O=1", 
@C0/SF+8*SD0>"M>72PQJP@,<]#-#_#D6B:>%YJW^N1  
@F?X-4+?!BAKPP'V,H)A"E[@KUZ..@B79?W%+49&.U5X 
@(7-[%/ZYF72UKAEHLHF_BR!' D<V#I(ZWUO&?<CCHKD 
@"CI+O]L=[H=DHI'A_]NDV[:JQ[@BN\86T* 'KXK)XB< 
@#'X:$R+C[FE#UVK]Y9H)UM_!G%M+W0B%D0O)=#.JTO@ 
@A9Y9IP5!0C%$HK;1([@2I9A\8H+;KG5['%M^*RE'#4< 
@1V70EFC@!9)A\OPAD*::ANJ7"#YL[?:PQ?K707:6\)X 
@'[DO1.8I&EN7+<'/.GA=5N0!A]A3!,S?)T6Q\L*+#9T 
@F)'1%I4CM7W*J!"_B5T.U_RS^H:GF_'VP\_S/SSZQQ\ 
@+K(3U[VLO7)W*=\NZFD%POOFR3EQ%"-O=S[W6-7?X4( 
@W&!G'^'0R27HY<!+OY(<PI"M)H00EM'(P$5WOO#N!7, 
@BYFVY3SD$?B7Y-J6@[3OZHY3!\+#-+H+_V+6#7)VQZ  
@R6Z/X;$=,O]<:)PZZ),Z_UN-MIY1VTRWO/P=="PF*$8 
@8%> 1+$[LY8'S4EJT1Z[)WJMH*OQ:R,>0#G^SE]Z)W0 
@-X<]\V;_IG3:C7,)DD??E5@8"IK:=O!__*2\;_R!39  
@,BV,H)N!F]X6S+Y+FY743^.!U5UU[PXM5_+Q\C+O#\( 
@3V).+UKUBC_+)$0&:!S7,8'Y1DR%8H'_#A_&B'._K&L 
@M(?/*-137&]U8%^7=CZVFPNI<,5N.]7B6PI9-GI5HA, 
@1IV11A[4TCI#16#^ Q@0U AI,M"1@(OK6K<+!3'$4Q0 
@BT^.88GRAT+VE@YJM$ W[M,*S9VF"=6G-<!LNA5<:R, 
@/Z-O<D0EAO0)DF*2"W1.XX-N0&:.IT,H7+J3T:U?8OH 
@,,4779K#W*F69:#51+66$PZ#KM\5/$:5"+(=P;!^9E8 
@<K XWSJT@0[6F]%.^N?[ /L,.(/R! ];%X1UYH+$N^, 
@RIB+(>E 9Z23./'8$V%CYN#W_(/R\9L0GE2-J<_S9N$ 
@6$5JUBF[<@_B"#'8OP1UG90?WK!5*K>L&2NWS>NR%]T 
@'Q6YE5Q6XA @0-?+8,TDCHU2PK$L\T\<<L5'.XRSM(D 
@(MJ [(2R!,#]BM<T4,.KL@YC3CM4(7D]1!T>>';-7]8 
@/%2GIK[K]%/8W'0]Z6@\,409,PIC-S49%!((5@,.$:, 
@-P.%=_L9AUU1L%$;]=IE0BL.]RB-.]9;#&?0P$?YRKH 
@PO]-2>9OXI0DLKNP^8%-G)MHQN64ZD?LQF9-W]1_0C@ 
@U&?AN-&DO+PK570?"0O.SZN8@P%,K^P8TIZOA:S_]N( 
@,G +J7  OWT>;7O/B:-&P&/%S*,9EA5JD H,+GS_,@, 
@LI[N_Y'?@KJIC=225NT/ :F)1KKU\1,0[XTA8NB*1%< 
@"-I]]MM<?:K%T$<S<'XI+D(&5;ZT7"0?U@"B, Q27($ 
@'1NZ)*HD8HPN1J"VC'>G 8WQ4"9T9B.).*Z!/XY)IL4 
@+[&70F82+RPQE_1 :I3FH%EJA,(HS4+!,4!3-T.^ 0< 
@Z+S4()G:JDA>=:#(N>5JJ'7:4_8/GY-,TGN^4PM(:\@ 
@-8#;*QO2,D$O3]OM5L>RI%#Z/18:H!FV<]MZN!>,A50 
@>+\1AJ[F(:U$FL4_?+1U:L9Y<P'(?F<)&F15K/P(608 
@!7KA*OI9_X^Q<7T1AFT' ZE3U(RV-G:C"7?96]Z"X1< 
@X02X39HXL^"'$S=[X1D J)00OH;I4<U$C=:[M?9ND@  
@79'W[M##E1H0P1#8.6N8!*'+/*M)ZJ9$+8O$J1'38F  
@DKE*&AA"4%%R 4M,>0'/O_3I*?AZE.3)C"]G*;LQ+Q4 
@6$@@#;(5;3G1V,!(C?T\H:>-<\[C2[SL75.VR>;JPV, 
@B(?/,? K?=$1YZPP5/*PU<I+]L^$APUMEB;]98!7D;8 
@GR2F3V>HS/K3E57A=1"8XGU.-'K&?Z"-];.?>(Z?(2@ 
@*W69L:9DJFX5]#I'\AQ#__LS?&.C[LL+IE<R$Z]]L78 
@OR!A;.(_\OFM>MM:3OQ8A-.T47J$V_I=(^@+ PBMK.( 
@+::RZJ1>OM=6X,MA_$ 0.>Q8N-X/$<)',O=]G<BX-J\ 
@R/7J,&+Z4P!X V;^55TOT\RH)!F=5E"X@_<,SMV*D.< 
@CQEF@ZZC->6CN(K))&#'=Q"4AZQL\]70QQ'S\2SEO,< 
@FEL8]V5W*3N;C%E9>W%2Z*RV8+M+B7K+GWLYNW%)+!4 
@^SRY@J\FX=4*UD'UE\T5U@'E-]";(;YH;%J#TL-Y'?P 
@)IB9>F[*>5&4OG%>]*P-.-SW9QP!WZ,DF#-SS=2VDLP 
@:Z 2!]"G@>&R RLY&0DY!?ER'<-ZQ7F1I26C$Y:.#UX 
@_+=?]=4U_O--8,L4U6+_*@C AB[R7O<Z:MWX:WVZ3(T 
@@W^G#9H0[\0[TH*N#VH,^OWPQMLXN(Q4^>BA96\_DB@ 
@88J?RX4^L',W<>#M:U#@)>]PLCC!T//!6UC-0_VH0?D 
@4W=EUF,\5HQ&/TE2>0+B!?DUKQY*1$Y[>RIUHW?U6D$ 
@*]GCB!!HN%,K;J.K0_3J]J(L@"4!!O+#<V_I6B MK!H 
@C&3[N'O ,*UC6&Z:(RD+[<I+.AV]#FEL]XSQ08<.P@4 
@$RUM^&WV&DR"+%J_& 1F#>%S*B KQ^W@^18V+^ >B!\ 
@6,'K<;<$?.TZF\&=VL,]K@S&9H0+HI( !&L)F^8*;M  
@<F_@:$D&XV%>O3]A*^0 B)YDQE.+('09!,*T5?-.SE4 
@_"B+QO78(UC8]QA E0DM)@U';]N;7.O4]*M&<2KJJ$, 
@Z70)QM4+W0A0Y;:RBP1L]1$:2)?@0PZ=2&G=+BY-<\$ 
@C2'PG0J#9)<A2AE @6U3]V][ N[$;+$2:#SQ]',#6$\ 
@+<Y35"?S:T6PI46PD5YR%H>E^?O75/%_[SH\9)V[EL  
@QV![ZTP@FGV!3Y.1GU.)E>"!>#>=QG3>CAIL2X7UU$$ 
@E"7N@1TO;XYBT<2B[./7#S4@;456[#?1OOKB(XRBH&H 
@L7$U,KEB.(X_Y5BO^$DOZJ_<D<J/X!&0=!0\>#G-KUP 
@=MJL7R;^3/% \056JP$+U?LV.J\)A?Y.M5M]6JHP;BX 
@ )O(IH0ZQ))XTE68B,#]3=B3=WD(56C)F-SX& +0IU\ 
@:M*R>C)6>Z"DZ/"<[8QS51.0P4!)>.YXF,ZPLN,%*@H 
@IPDL^4\*)R7\'4\MX)+3>44I DP=OP]!9G>5=K5PWX, 
@.*><D^816VUWA5F([>9#=>UF C\'AH'!ZB?T\-Y()ED 
@5[(;9-Z4&C6BII]_@7B!65LH]I6BE%XAW\/K-/MDPZ4 
@QN0A?IE2FSU%_)0X]&B-95!N]R1C7;*LO1M$259$K@\ 
@II_]^_*ESOPY*.\.G.R1H'4G5VAVP[TG K9I>1?G0Q  
@RU]B\EN?[=C0EY1"]V"9W>D//-1'3=<6(^ 84YYS[QX 
@9TA3<DA /=) NNSZX/\0.H;4'_V@;"C?ZT3T0MT%^S0 
@%C\#QDNAT/K;OQGVEQ(!U=+)C-_1(0?C#\O9G2C0_N8 
@ ?]16;TN,2=NC;NCW^./::QMUJ_G7# V8Z1(/ZRB.NT 
0,!/5L'/.0>KAGN'U2J6Q#0  
`pragma protect end_protected
