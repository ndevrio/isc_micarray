-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
GDJMItf4vIVUV3frvV/vPIKW/wFqYg2BZVphC/2ybO8BFDq3mVmBaoz1B5xqQunl
w/yiyl62gxyt2xGLe11CaGf7tOiXPOvWIAE2EumGGpn9iJUEFDUWEa0wAF9jVstx
ZrJGBfsVBSF5wkB1LbxEWswNdjJurKD+M5sTGY2cGTw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5088)
`protect data_block
cqyNxBdgJ8amFh55X+JHlFVMy92Q7zauthZMze/opkAZn3Q475pB1f+dnMcCJRun
D07s+aLOVTBOjZKYLJGFnNmtFxdWv39aFcE8jGzHjLdqqTSIyPmGKBlV3aETyib3
hpz8oSUctVOGhXkW1bmTivbDPRt9UXn0cfB5RZo/u3qO9rqP1gWE9vEUoqT7aOPK
90Za4kyLhkgDpDBqu+jEEQ+Zvb4rehigTdBY0wY7a2nP2jBtJqMGecaRAe0DMdL0
ElJxENklTOYL8rjC8o2CatnHRNv9yBXRYhQKz6jL25K1y5Hg1X4wtvdEPtdTyjdu
s9aVOHZiaAeG0TgMYH8Rs4A+uAdr35Cp5YmvgBsebjmqu0iB4nm+1csXLM33FksO
Y7tn8jxRoxZ+1IwpQfgvUpf/UEG0xZWuauoJf+rexLEfDmFtustVp6lNN0mwvL2k
ZU8+YC5G38eWcd+S9Qk88/J9jyhGSuv1vhuoATPlwM+dxZf7OrRybP/XCnkFWjaN
DjkHH/FLcOZ3H17Oh309B+uKYZ3xqnicOz+uHfCQRd8eBpp4gPzLoEgQKx4gMOKG
ZAOTTBWQhCjOn0hDnQrir6o5q5J1RWRKLswx7r0cMrgwfJC0ZuZqSXBk6zABXAhl
5DUKPscNX0b/lacA4NuAmW1yQFzkAc9TZlX0aRUDM9P+AeAEgoJLJAU/kwOjT5nV
m/qTwHkqFdmSMUrOuDxWae4a27ATv7nFymtt3j8pb4TL4iL/fNUUulkjA6RoVvaw
Fs0/3JNh3Ja8+4TtVyBOz5he0klzHx1CaTolGl4bo1iMLutXrm4HvbnQ6TkvlJdM
q8NuR0c8znNAixdpUlRIjglmVszwyCMOP0pv5RmT2XEM8joGjPtqcKPoz+iLc6Ks
vFkrbMLNVoVhJc/+TJhs3/5cgGeT4qZt/LCZSS/XXqxEVyhwpJReU3BNYEcfKpdt
eVqL6E5gM4jCYiNjD1L75KxBvMk843VM62T6mYQjrPZo0DbgFYdKzwWTK+CHo3th
Nr9fVByRBdPCKpKLfArj/Xv/7EhN5uaCdS0nAghtVEcKzAAmqJ0EWxAHXlJHVlQG
e4riawk3NT1s3oO2SfCFpPfl5E91eSF6Yb8azo5hr0BX9WSs+0qbncaF+FvdWn2P
5EfATNRvg6nNnDfliV7XV2akNwMyMvSrBh3wgL8Baj0H89Gl0Dxinganc3MgPsVA
mB1KJH4ZtxVilxCgFFFSbj3rzDRsnnDlGRKfRh6ATlGIYpjtn3yIj5OfMavJO8Zc
dchKqc8icqwlwaNW2KCIS8KCZi0Pr4bSxl9PSGHDYVALX4NS9JvrbXlW1Tm4mKrb
YHlOknWKfpHA5NoPPBqWDLyIqztApfkF9nYmovEujWQGlIAlGzTCCeiKfK7OLfK6
jo9oa6Q+0RyBaCyCFRdpUpugFIVHjFS1Rnz9J0rcfw3EtbvzJKGn17zOi2upm8BU
FI8gQhUkB1H0zKAWs4zlwBfxRPftYQH4aqpdn3os66UHgi1LSNtrzephSiYg9BgE
QxicrPG8Zjfci2WP/21G0jYSBLPqtn1CSE/HiO/wCd8Liipy9Iq4QnWcR6BeKZ1t
KPDtKO5EyRxNQWp840zwfuCCwTVJU6sVWdp8k89ismCbDzqeF+cZrE72xAxEEeMe
6K1Ypv03j8++YS1GfuwIRi9Kv4j5KB22zOCYGakDr9EOpUiAviTspDlMzLDnx8U9
Vp/hqapRoIB01TdHXzDNxto9gowW2awQmYkwSgCi05GUCCXjLraCWZPVNxBjRcyN
zbpB3HhlApo+ZGZ7jR90JxdPH2dLaDaD0cyGsMZzPXSoNLDgsRCwTX9VFQfthcOU
7Qn9PFwo5uS7lMp5p4jICoO+pJwwFK/XKL6jiqaT9P1PVKcF+LxJ88IZ27KV/aYu
euyYcXfYGfsZPVNHKHTMB8Dvel27HVLa5bkVFs4X5bsJKdqi4La/6a76ySpjPckP
p7XcvBN+fbihtxoR80r+v72k0o4V44YjJeBgg34B55BI6iHsK31fDm58vZfHR2zB
mo/AnJLd8PdBRx4sGFVDrToJwIzHsVsJr4PS0gwRlYsHvOClBLabVXghSUm3eSJD
HKHwkwarWr3fSbY39ihGl5s0v5gBK4XG7tbUbLyW+NBGsMK8Bw1VYy/bLvTwCGzx
rCNF41QdT9n/g7ra0L0sDVzEA6aiaTV0ygjxQLub56F35QZPD/ZPPOpVD0PNxD4r
BvnuLLrQm173pEv+uY5m6sU3wfBPOEO5HXtfQXrMOZ+haLrLNBBJMOdkrn/MN8VK
vWGBH7j7sVuMKNfwergI6jQnYVsZJrDhR7IXK3/aPQhbYVyM66xp0dR9QKLWHp2e
49ywj1501l/TZpX/M6O+0EAswAo9LCb4VVXCdMKJXgi/CSttk+S/64rTylMuDHjN
DvRuTt8aFhYLc6R/wtIpH4b7Od+DcSLjrBptNKWlASvJsUeiwCCuYkTetd6c6nGc
5/BeHCcXK8aZUa4WPzi3uB56R3wOVlrolD+jtXYch7IupF/woh5VuRDfvhuf+dEy
v424G5wjifXARAPmHwiCMCv/ihz19E+bX4CCQhR9tUVF+QGg8mc13S5ntQc0Qv29
Njq5qJeEpMQWOltgcC5rLRN9B0nCdnkmPVnZOhYA5oXkXnuGNQzDvyWzlhIiU1r4
JeiKRRK2IWO5WT8B3v6wvLkjOvvNQs76ZjnRH5vItDJ2xcE0zTr+1IeQTo/eThh2
ik0bEaC2s559vHNG0zMS2fzJxa6cxsIkMRbE2G0kiR6jLuTZNbOVSZjSGFsRFHvP
LhDUCP/OthD6GCnuhPETbRAg+R7gzRTTaBJPUUvkMQRQ8O1+YALkYKklBv5oT0Vq
Z8N92ldiEoM1kag2XUtnio0t1FPh/xHV8/3t7JAM2cTCgBlqy9BVG2bOXTYBhsaM
Q1pjXEoDnSiDyB0dBnnwujtYjx5REaOHPR+/b0CffpaD+bJ+j86h64e0bJwIqncv
QlLLINYWscEnFKVAjemzKTCIEkcIKmNZVh2R3ALIifCWv52uIUSzAjZZzXkfj89j
KhkIb5VFvGI8ZTMNpQds7j5ThGbOxJl02eJ/X1v/k4ASaJZjXd2j5JZggCI6VBlD
ZJDCtNXuNIxGyGgSLT578cvgN/N+XZ/+5g+a6R0HN3XUKPaX4Ok+vdzi/5on/EQK
aItQ1GOHmrDwC7PopFoJY/kaLu+jxiX1Iygdat/do+bw1nuOC9lUzPadGNSg5cTY
PtX1WoW7dQeWG86FfKNETb1msYLhwu2mEI46C7OytHzk77w3IvAJ4QwliIR1l3wL
lGGbfbUcROQf/kwfMp0jpg0G6ZC11G+VJnPeRXt57PSEtJ21Sll1oKQibRetkN4c
iVcBYf3wmSePKrmOkC3pdeBdzctGL54LUeU0wuQT2NfjfZRXjKpwXzxcxKxoEnkK
aIsdxCgxQRTfMPfMa9xA+WvFyyfCKTYT593Z5vCR/Bu0S/opVqG66OCOxHsa5ogS
e1lRyMZSTHXJAaKnO3T02pI4XP901fnd4sgvFtcAN5pjIXZsvI5JKppMM3Z9aU1j
udlCzmPfYXVLW/GUnohPQT97SYFvePV+IsdU75SNo88gF144G1Ng4i7Bedtf9Pep
1AGINQXKrnmBDESeJ3jKfQRhLYagazC1lOSeYwuGi6UCYb2Zo5yJtnU7C3bxcgAv
wY35rNL/VvTVST4QKs7lQEKIYRbFeJ2SHYQ2yNEn80etT8EjB2C1J25VtJPgqr+k
6fzWwCBMtOtsmFNsp+wBh/b+XNvVr9P4Q6ycS7qTVehk/inYPsA93wg2SJMtgCgq
ADhyB17znMkdY6ZymUUBEbpPHB3lV+jYcbjAOvBIBjPju3GGVLLIyg63eG3301wt
AcMnKAJe4FVScPhADhfKvT7U80O2whUJR5pg0LBM51hGF2FaMWKdlL1b5KPj45o/
xOfAynnhwknQ0awCxfNk4iBAnZWuEe0nPzplxx9wQUFfbSzGImyCryjZB6E/FdWi
LdhC2ceAhf6RZ+oTUWqbz7jT1qWXGAPbTaZlSU8wX6jKK1TpYRKL4uZtGRJR99rP
/9Y+fslbIPbTZDWvXpG3QBYJNDbVMJCimOg59qnpsSCOsDdNImInLAj+q3uBw9c2
YTmsKBYfJtJsx7HA04zO4dN23iRdSZeRgp4ZxlMvDSt7BZ0aCvQM81+jgJTnL5AA
jLq9J8gRxbHUm6CvnplIyHLEPVpaVPUnueR0rSARkT7Y2XLhBcFOxakmjA8Sb6Xq
g47Dep8C5Xs5SrSn8igMLJ7l52nTVE60MiI0HwOZEDztYbhmaD2lIb2a8ekXah0k
F6RLey69bEawsmSOuGDaYPY50K5N3d1bt23e009EF5+RcYIISb9EKhQuyAPwelYx
hodHdKiA5E3xs/+2F3d6Aq4KSB7/w2+t3S5GIjbulNKhgRB7MrfCcwqp6zX4Vkjd
4UjHZJTQOm6JqvTfy+yHzW5SOKyK43NX2MU2DPW7Syzz3lKhL7i7MibkqD9hGRW2
kfWaqaLWv0v7XO30fHX1SWH6WSnGGVoNgYZddc6LDTY25ATPCrz6vzhjefuDw2oS
3XCwQTxleGtnwXuyPx3UbnxjHbUOqvVoflorAQvnadc10EAKIWRIb5UXDwn69bVL
OonCj1mpIzI15b1d6cgGUFxZg07UgjeW/BrvbUPU7sR48rPav8bW6/86PwkhGDBC
/Yk3VnEulTo4bPkStB6Xj320Rrq2ex30Tj85Gsuh70I2REFuASIw0qlPTI7aOssX
+nWAIfFZn0opgscPvO7PeH3EuFhINLvfhyLCBS0dOIsuIEtugp9BwD75TSLZJuFc
tfPpt0DdGMPk/F2cIF9Vi+X3uTTvcOo2rbXSlxeHuzZdyT4PR4+9sym+wHlhD4Zx
Icn8V6VPFXt1JyafkupB3PApblQ304M0pTi+9T+Nr9xSF0vWDpKQD0IRKxOrweKr
ENTGfS7/PR73OwphENZVeMIdPALDjdEzsoR8auvNR4hBUxmiemtOtp0BQYS8OTLy
UZibOz/vwOEwNZQzhDdDKD4WIsyGqYryrTkhu2YhsbEmkwNYSsMmEZJcQZyQdgNH
QdjpHpv7NqfsCXN1qgK4wvl4EYsRhFtB0iag6DJjAkmLAWlWX3cWBmtGXYelYC3H
KyEQ0cY8IPSPSaV/rKEbB5oS9Cp2eIBLbg767XhXFZccTzsXxAd1Lh/qnyzGZ47C
nGzGPrIihsDMC7GSYnC4LHJtyfUoL9C2bgsTYwMCY8s9Sct/CmZHHS4hJcLUTZFS
TT6fjIukk1FoPgB7AdNehLB/rT8XNj4Qe6NYAbAxJyOEhxWbHr1TXcu4usqRphbb
OMkCcF+c2ZCihtrNvtdvxVlVGwJxubfRBgiX1YMELPGTV8pGrLlXdDaBzXOjMRx3
Tr7lYdhJuPxSoaIpM8z+M38ooUsn7MI/2XBgOqy/Q9tons4LfKREuHoZGIW8Uuri
Er/2jNxoZZt6AUMLV17m7QbGTCmUALpPekI3nMdPYHpdYR2hdRdBSXpgYDlM4GBW
Rckz9mBohHAZxJxAHm7ulT3hT3qgwrHui4rsuF0PIqEXgrqqeXYuJ2Hl6Og5LwKk
hJ+M6Rq/uVWV2v8dI+J0I0DtMyhFM6TrDHjiRhosNDjBi2akVKy8YC0vlFNcV3so
IfqQbJEfuRWs6jNJLO5ShYlN6IHjIoR27eCJZE+9UQPhHKFEaNtd8Mlr/lhqsQfY
EHmevzpvJarprKi9urgyImCIh7YjRroQfGSqg6iPhD6JhRN6WRcnAd6wLtBqaacy
pZL3t3lScU7Lwx9oE1hTXRe2pTsB4tm0/SauGNMFRWRVmi4CNU/6WysHSrUrZVI/
iLLzdEOchClweZpQSOa0eR68XViRe3U2MOJOG/7UaRPu+A9MAZ+JSUFD0LMlRqqi
srl631owePpxqLlrxS1dA+XLidqGzmvS1xiEcKUh8AtRd/g6tBpBkp6Z6LOWJQsj
HwkLRD6gy++pC8OgUdyjbNRxvMAwuokWNk69caQfGnQ1fp4o/uS1Apjy92pTbC7Q
UpLy1832YiacrU2sUeRT/MtcE5EabVY53eQbsppngV8Ck5Id2GGmqisweyjYzE2A
AAIIGhtaNAqqFBHbodQYoZ/kKSfaBtj/qRSepPXpLA6udtgczZ0pmwjsJZV1tInV
ubA8UVtLJbe3Q3atXCeW/8RN/d3WnQpJBenXmBsr4HWrMojTOuzx6OEhLZGi4/p6
CezCVjHw/HUMAs4zCdONZj9CGxsYcuCuhMlcCc7ctgh48EUOj+PvRa+o0iazP3Mf
HkQo/8dLs2Ip16tXHD7gpD6xHek98wCeNStKIPGHxY8LURdmx2EwTIGC9+lhxhpj
t6R1+HXqR+yEVhPrJ93VDBAslb6IGLCAYhxILRJ4yOfCE0eVeNcAKgw3lt6G0ffG
QuP4ma+tk776XrFktHKBUdNFJvPLz+CVk/dQpFnAUFhb9mJ9CC2AVGi5HufxGTE/
qezGYpszBQiWBExDLy6QzQvYy1x+GxCK3uqDSFEKUiqLgaWiehlGyRmQ2415oy6O
8IzNaiPEl18n/WQunO2JHe61ajaF8AI0vU+vWohF9uz24gt/hY2aNtwj6h9E2tgg
L3TraqXvHnyYE4dwn0T4w/vV4M908G0G4ctYHYQ89AnGK8LiNapN8C7HSwijwTlQ
T/RkQYAGdmFBWMFcwXS0n1gbyrBZRfFZEIELxzheq6wdoRcwbrQCVGNPnmFXJQ4d
`protect end_protected
