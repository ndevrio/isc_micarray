-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
PZdz+uNG3fydKTkBkppQ/YAVjBV8qIyDg5TbbNsMb7QfqApafHgblMSPJ3tMelTYxrWmGdNYrjck
XbrlXP/ZxMXZCGgikwlshRdj+aVNNWyKtdUgVhjYCdoVpuIApZlt8K6Fo4yYXxdn6fICM60UluHa
d6MEkfTMC5oGeGZUB0yv1NCX41pVERZo8b48AvYEmqPlXsv46d+ostdGK8sH57GQctJsKHPWDfe4
fT7wxPHH4MQK98+FOzIEdGPUAUKyQbXX7oNt8ZgEul5V0CJOzt+jPd+9bbq3PJQ0ZtOuc/QIInKa
wSfWwVwMEMLIizJQ5XV5kMuqc4Y71LSLv6f3Ng==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7488)
`protect data_block
at+RwiecccmYDR+kYX+gEfb205Hp95sn+nWDSsRjkD7xW4YpqQkHfQeqKnzI0T5Hv82JHHJEqICi
8CwxODTfSGYjL2nk9WQ2dtLqgSASUo5eh/GIsigZmb1T9cVoWFfRmfwIGgSU6qHpLNEaaqz8rhbM
pGVWVvALd1UezcWeFj9pK5ARLVkuHTJoBFac5WQJKhHhqgQuWST/n9lBm3Ms/CXrN9JRSDDuvVsz
3sWlvPM85fhN5SY4zuZCsDBq6HbsOm88/G6MIigrdxdCQIHbNS38j68xcOVHrabcASDmsjpnMlrh
vyY+P/QvH6UXi7BAmeiDA5kXBchRJb9uEXWGpLJBj0bRnjkHpZqmM5Qd+hyHB2mnUNb0UJV9ymN+
IokurLZhB8fQYJAdtLFmMDrGFxb+ySCvSSiO1MyOxJ1qtdGLP3XNp3BME7VkgSQEjcn+Obnn0o4A
nx1Q88wNua17Aqpua64g8i0+aCjjIRdWwEEoDz05bp9V3ZN0Z3cBNZWawOctFCjcIN/hDsS2J9m7
1kJBGBpEeM7u32Rw/BAxSNemDdinq8HHRmwpdhOi+80ZDwkKr5qNHs+diZ882DCEXnwy8ue5VhFG
PqRVf5el5dvP++U1SDW2nRjmb4lNq0hnGT/jY0sjpewrTne3zxH0jkeJe5fdslCaE82gE5kzkFsP
JIuuZO2KUvoG4zrckA1Hp2efOE7SLUfN3OHf3b/Byvb1QTQKZ+rDWd5D8kChXEqLBMmtRm5WqIUA
BVggkGHFUgFe0vwMEQVFdUQGiQPDY4EKU5KDSMl0iDSSwC6u1wBM32XzN8P2uKwLRHSgbyWecN7m
utrTCmuXt0IsZk6lOGpiMCduNEIEePTNxQtMU6p+mrH2/HLhE6RpUPItIAEJIxMFEPuIUfFvzOy7
suucn+P6E+5mdqbWfarZ12OYaFYRZYj5Rq1tIUnLATBx7OKTcMd+orTmuD0IpRhMKYIz4RIR9ZsK
yOawrzxsVbEDMLVnrB2u4QmQxJS3NohTwzHg/C8o6zqGqjqsK8sDx1E6bFNXzZRMta2D6bwWKCbg
+TO/gc46wv2J4TxzDCdyIZMJN3LtU7zXnjjaLv3swafDyMoxywPDEViuIjg/AzETEv2L3mVtWswV
4JTB0KDgLCz/IXSCgBkaRcRavoV0HuU+sVkLPfg7Ch36r9PIFhFWG+mOvvXhJvshhqr9x205Uih5
IV/4I2IUhr12oGA622immjslLnCaCJASNBMAZMN4uDhdvpZwka2BC7o/sIlDGr8nYa/SahYdn8Aq
yrJ82DLTiqsspe1SJH6YJV+Sa5vExopyf9fRj1zXJ5Kie2bucruB3PqhMm1jSJAf5PGfR+fzCpH/
tmXcz/ticTNzjGcM4BP7CMqHJKJxu0ligcj1GQuemw89Vlt1cZcbB7ESIVnpJ7K6r7PGP7z6lHZo
iTmN+wElVknOW8iRPo/KXeYHaCrRQxzxIoF9DEuLb12h/cqX+7CdESlNJAE3f9ODEqTiJy1zhuiV
gKBCgb2CWOags7FcXfxtE0r9BMNYnDJc0Ug+hK+ldgI+gL5XXW6yKV4I4nSjSTGn6JPoD79ytsDh
WcOVAEWqjPqDyS8y2439g0AQRSPAQxuigFZaYTvjRmAQ1zcpLXJYWWv5oieGnATIMydnX9sM57tE
CM48eoom2GaDC58y1+y1psiSmJmyspGUKYJujDgXKtcha3rS3JVRL5i62HwarYgVfWfConml7Str
LpHEi+/kdgJeDAzoEeEBzoVBRUYpSQuIhfb6KrjE+qTs+hvu0rSK3+kIqxEpfyb+x/7ejPKJK5xt
0caTfpKqxG5T8S4nVPkyWurEwfsXplVIYK5hMJElscPQnqeokSvPDV4PpGQvh1I8W+GmNyv10/KD
jFjvJc+H2Jin1IHHR5w85VtErbSUEd88TXBkReNkoMl976MVqDqsk67QCIB0oAc/kg+8C8vrTO79
OHTiatBXGXyhN2xrK9I9QSeCYwo7mDfII3I+AgEqAMcdHypN5Jw4UlKCmwrt4cWcTf59W1WQjaJg
vr6uRQFUOqth3cS9AJR22GeGU+Mc5/brSx13HErPzd56ZVvwjTV2yU8QomhvpupMq+GGcZ5/bKjx
R0c74qp+z+0VvjzlhzmpIa4B76eBCg3iUAvvlA57nNar6Dpu+ATvaJsJeZTNBOtaBUhvREc7A+PU
ZFjpOTL5SsNjwnG4bnnSo063sli00T7ypnVkHVd4duWz3ViGLQN3ZM5X74p5pvMDi+yrZoi2s+9k
URCnEi+lKG9WCUbh0RU5/BkewH2jEzFJ5u7VAIXwxVij8Ur4GI+6fGffeUYUUO9NnP+p9VkZLoPP
SYcJx7vaU3RsQyptwsekd+gSq69uRzpT2VBLsTqRiowRQcFx8WtnuZBy8rcCrGIddc/Rbv7bDZgV
ZXAQlxnb1bt8lQWSbazH2PcsrNeCMMLnhBFdAtFICBgqQtNA1ugGnOzun1kS/0ltgj48y4pabZpP
5SEYk4QqAMe7QSsD+3999QPoVJwoPqzJSUhMTz1mayBeSfb4DtIqGw1siDqbEkypoBOmlCmW+WTO
JG/IrJ/PALTD8RG7IaoLzPJxm5YJ6R4Erqr+9HZVNLlpdnt1MKD1ZgGiSKRtZ+ILHKzkbQcYR1L1
1mM/7MQM0vfc/3Cm1wk6sCL8TRwt9bIRCXGjO9ZNpeASKz29ubLrkj1d/0ldw2amaO2NAXzxpwJj
cRMrB9yqwyH2YUMof/4hJtLOjfEH12GYhlrjOnq24INfE/aD3SjuOE8R+cRGrZsT/kfcf7z8iWl5
WJex/IfMrQtpewFzZt193XW+PI9uRxNq2xAuKufwaBqzDJbCo/rSl5s0MTXYFVeh3IJgOi+/1tI9
pVARSOe7vlm0wrsx52cNmHQEDY/Nq1L7ssDys2ipecdKJifdhZzu/to2a+gAWuuzW2wSVgCpRRJL
4iF8FDBkQvFkgn/d+gh2PeWh+9BBXd5qGEvULfupQWoNoGR+rMYOTT6azrOtgwYdBacmPgwbaho2
5t0w85k92VOJzfwICaFcmlfq7uSoRnsZ5pHZTsTIM0Qg3subPMOURUJyVJb1w3dfwS0mwVdqmzWC
o0r67PfGSHZdlp1fBzTH0S8FLwT6HumTLmHh35QfcljosHTPGYwGSlKOetELPRJYK1XG/f84bkW/
0jFgOVK55lJQsYnkj7/2CY2fAH3XRaNvMLd7H+BxonelaAxCFkyA3OG71F7DPE19MeYCcIkQ8Ih/
Ce+qg7vtwCBz+/krNBVQKHsnVzFJWMvZnXWJIxEeGBlTETznHqdJuU9Dq9OtuOr61u0RdDWCTmNj
GOs0XGL8weuEyUjQ/kTyMMRnHbXG7sD3uyalOw96+tIclQdLcQFmSDgqce3h1/EDZa7fruDg9gAZ
TPZU+PWBxbO4IV/LEyuabKNnP4OWQUBYNgJjKNq1xQgiis00OSf3XaUHR4KHDqfBGf5CgfvgDF5j
zpYFtsuNgEuWwWDcCbNU0YVuW6N/eD0nvmpBTbVFXKgQvhjxOoDSUsNUHeaIeWMHSTV/ZJv8m7nl
vtqF4FmIJn5Gld0yAPn3OUENLEQU2Rfh+A2Uwu5DI+WzNImjKx1V+zsbxm5IuFbespn+ov03TDH1
x5ObA5BdYN9//LT2B1sq20DhUsTMxijY+OdkSJmsUViGUB3b5IL4iktcikfNcCSLSH+TTh/8IWQH
b4M61woXAHVx1Z9ia67Ym8PZjHSuO9mFa44OMkvywodKSVccq6OeFJGXV0T1AfXBF7YICKovNNxV
I2o997skMlN/uroObfTlYLltjxqzKXb0j0nuKQRoBSLfvMMEHLXQNKqD2ex6bv+AaEMi3BcQ6o2j
TX3l89SX3m44y9XY5famO+3sMCZAiAJP3GHPdIuNGZYbyZMLe55reFFIxeQC7LVo22t5dnurY+Y3
O2i49XhbPBlcUJBeFKssVi9WOjWxL5/HkcI7BxfrIf28xrfkqXJvRlOz0rV77OPBgfqPh9IOZUTF
6amWFRpqR5ZUFFSiOqf+hDeBRQ61f65Omfq5oVT/nTjqZotU+bQYCuTK2zJ3A0aWmaiqR0ex8FdS
kwTJDeQSQyxY5eysK/4Zm436qElOxy4tYNf2WXf9FL25QaCK8OeVJq4Rvj2Is2+16eVOUmtbfybv
Tp+WNm4F68hxu7nMsESbs01oVaJ0Oi7iY7GDiAThgUoa+M1GoSGSRCcuA7E2S6JetkRgEMSKtpS4
05dUkMpfi+M19rNrHL+cr2dOWW2SOlnydOaPkxSNZ6cEcB9RWdqALiJ9CObmneCx+GZKFg/AO4NM
QJNdRS48n5osk3UIyaP17kAlILRMSlTzlsLU7Hbi6wPgLu4u6ffL1j57JPh4hPbcIRuFYLbw3HdL
dhMVJNRArGZEj9YFRm/mYSLYnDoU0jCB4Nanc4xn32CefhV6b6K13EOhQ2EWJjJXGsbRfuctDfVn
ovI4geV3XxAjgAssZ5skYuUrDz2Njgk07L1eWSsXWAgU5YZDgHEfKMJmHY+ggHdpR3nBjfnqqmaZ
YirTNRNw2kX+25tigMJbZRGPI0pRRr7rJz6yfcFWxJIZU49YE9FWYuSNiz/eUFz4myJMP2wKQ0Od
TgAAWY17Pc27j1AGVu2uAJn7omxP71fLwYKFUGmbW4g519vgfmRQLmrOTd6awHOB0wXjJmo/TWB6
XGV3/VM1ZTcw/4YnmAGvEUsyk2LoICr6cmu7eu7p/V04ZHY7EREnGFYAngF1CyA9oesDlPtsct9w
eduHnsjrZ4a09sKRVTByyXKm5emDQgne/J2kafvA8Xy05tL4Zm2Za2MiAK110eKBYyxdpvLNSlRS
2qvMLgr06cW7RjclRvSYaGqJuCejVFt5c2P5LG5NL/XjNNqcktxh6zeIGxmzyOElb0D/19/QZnUL
FxGXpx+0mGEd3JnpnDZt5GFFMAXpU9OmvNabyoV8q404FU+BODv1qUg7QtzhCo82j3wGZ2PHh6di
TXJfYFs84smbIrOZwwU9ITAgjR8SWLV5QxmAVXMzItny02KARYdrRSuDjvDEHHp6TEf0nai7Nucf
0qjULWdRiJijgFng2t2qFlEqu00nEQKxAjIu3WwL6wr3h+V8wyAnAfY9nOCwuS1QrfEhPDXCUuQb
P+sFphq3DWe6OzY1dl3Ayv/eKPLyq4gedEtaFrUwhO42C+Hgjy5U81TVWEdXt7LTojrEKiDDy7uG
Pfp/y+xzuKAtRCBsCdWWTGp/irV2lYkTT9Z9inEuHFyCvko9WGm+YtgoVLhwyAJb99jJvjWkKME5
R7YnmCZ657P7G6apKU2J8BxHAig0EmW+cg4cG8sKnEA/1U7IgEScWSknqOr6DY3Rs6QajpxtvdnM
SFyuIzFlwmBPDlqSHFVDgsCNj5vya1RKZilDpit97K6C/W9QOBrDYdRCr7s2+RTNwl75yewJ9Ies
PftI6MiQZRg3TfawZMP2zLw9X8z0gsot5ZHA9NdQUr2PxIdg7S8kD8lUxEGD+g6a2LJWiCSEHV41
tLyDe7iwCmtk+X68y0FzmyEQ/8NcNq8+q4mcgY3oBHao/RO+XFl7U+Wt1wnx+1Ye45ZYSwj226Xp
Vo0M1ok2Zfej4lZjSBMkXJnUp5m9sFvtlqXGptHdBOMvRXJza0xrMWp5sDsSiBJUy1TYZAy6BwOO
3ENK6RvLJ4NmLvlpyqBdNPY26QdFNmxQOd0751i5AINn4CD3VcpQvivh0yOTI1u79JjwgwuCmSAX
TwFzmwJzqOhZJDyWOPP1DLsAuhUixdQqKCfAoj1Akp8SrCZ/KdIyJAq9cIHveaijDAjQZ506ptmt
qpOJQNqqrAp8wYNcCHFlPnHk+fHpDVzYZbgEZYMq5frFfakOsO3i9Gen+6pGTcaAsE51c2hbVKTx
f6h02cKJYsor21S91mHjtv/+Bxu03QveCz7iE6LplFIlBIVFpExH0uhxJLmc5AxQTfQsj2HVYYLj
RuCGpRiYtP9ZX5Izr13WgIhJLJhn/aXWZ57+5k3HKDQgGBHufNJ3XvgNeopOYTQaNKTI8i5/2Nuw
JVelCDEdmWIYf3y0uWSBaHzQNx297aqzUAhKPuriYs65Rv7B7J+QlNFg9pFKdHZLsg2pFKPr18zX
H/0UamnrEAUwlSP0syfL8aVi11fvFg9lZHTyrBLQfMapldZfuJio/QjbC9Zy069Oz9ZFTaZo3tef
q/Uce0A+lBuo6BPRbh/xyvYt2M2V77GbCffjwZ2aNAhMl1pA94LttqMV98esRNdFvBrFxGJVKRjY
crOH49ytJ+LHmThyXV9qzxS7GIXPvrpHPEanjjNa49XOkyqU6pWlJXNq2n3xA78E50ZdHhJT/gs/
/S26WuhdQeInTagNpsQE4fk1cqZG//fMwdVjf12/1OyGSXlAaeyDGbX0L6ELOYwKxVUgPMZKIG0n
3q6GvnroLy5ADJw6FyXMVSqcS55G/1F82bAf1GNJER5qB76ilgYASPbFCq5Bn3x+rGSKpOZMHxA1
jHF5ym7xozSV681DXwCLIli5Q3Djsz0fLFk3uSiP0SkfGP4XJQThptZVNguujeGpfVRiisqcpooD
ioZUf3z6N5OY98c0T3BeblAm+umoJXtFUNG/kRcgeK/F2bjtb8MFGHJKiOUvchwD0QA77yncP+8P
mU9F9EK2pS1rChaksSiG9acdYS5b7MeZ6inPAB2pbqCqq9/OkJ+uktH2o4HoGdhTejo6YKSJJxtT
jUuXgXoxHXqrxZd3wFPLvbp7R6zCi9YDQCj23BGE6enf/B5H7G0QoXDCvl4iJz2IkQgx1OTZWDmg
iQIezyYdPdoiu18t6Ij4yrGTRPUVyInlJ4nV/Hfsjc4sT+K+MhKe9ZXqM1h5ia+ekxfzOM9qjh7A
VU/S07k/6P7G+VouvO/iq5RGuoagxmkUBkomF5I1aWKneYYK1VavsmtGj9/don39FGesSC6ojtzU
+Y6UmvidsuRG9YEbz0wQCopvXIf3a5bhPzbV0M/iW1JH/tdGDqUD6RP1/Z8Qg8R82fWHMlMs4gwS
AuOttT4zkYI1gK9r5LGz8tK9NAlZL9RjAsP9+OAWnLN6RxA8d8Tee50yoNHQIYhWe5vLE0/xOwuc
0oxvMySwx2votv2tBDKtzON+OqnCqvsvaYAvxqat4Ru7161XWUkGKdXRBsdT1YPwFV35f4NnN9Cm
NYvsFU0iKXGsVRBfKrkUT9F7SpWDVskkAcMoAGHXacY94KKe94mwXFlvUI0lGHstQYr+oBxrnOAb
66YZPgVcndCO0PcQVgMJ9CdJJ3mh34Ripnjzh1KlFFQaSjXS3Qwop7rwXhlDjPkG/8MKS/AKWsrl
EoK820/nDfD9UU0IyFvPd6Y/H4gsx6oGKjG8Veu4u6AutboxRkQjfk0NkvdXrPayRb/+pRlicp8b
wrapJXkNcliSq51i8M3dNaTpunBnBPE8TR3WxNiT6fCz+9EodVUWEvBPQXeN+e4C3tdIcXxRgAMg
P0mcqQHFybkpVQuyOxrtfq/OpbwIv3vEIiI3+CQgx8TD0QWEvorFMo7IUhej5ZR4fG7o1oOZiKLm
KVyxB75UFAc5lw82feCQzY0uufHbI9cNBGRxMkSK8QClb+3H8K9lIl1IT8PJp19Cj+2u4nwyLTeO
7OPqSMBwVTuspKbVG/OLZI+5vQsVEi/CCI03V+l1Tn4yTsilmfxLdFpYb3yTwap2XbJyxbqRbDFx
Mwj9sECE5scTODYCI/IYli8FFq8Za1ed6qY/lH16vQTxIv4szrJRWBZjx0HIhtHQy4UJ9/qOdhwT
aABekimIej9mHM9HFo0GAt0GdkzhJxy3Q1yM0z0uuKkbmt8DU/NdvtRvmMLqqZ/EnuDQtEIeBjbg
oHztAfqfXx+6ZUsl02Q3GhQvbW+uX8qnHm5hQQVN9FMoa/yBGj05TdUa+VNKnagATJCoS1/OnrOs
4DXQw3OyJJctB3P8KXjse5rW5L6Ns2EB6kRj11QCTbiQakvWtBlFF2GLumo3zzjZfSCzErIhPpti
BDoTYe9h0ALZzNXylylzpHxyIkhULha/oCxOey9ckR2weNgaAxI0IobEOZMnUCS9WRxjDLFali9j
jed3JFWZ1EAapYZ6Duf41MrPne1+Z55c0G8Yd2Iz+YpgJ+ycm3f/yAf8vmKqW8daGpDQ+jaxxGQy
Ul4/bANDph83d2Xa6S6wfVZWY2W9I2qOncA8osHuMXN3lkeddJRJ81o6H5sdmSwmMSycg16B+ciO
KaBgWaxuMvURO2APC1PU8M3NjGmb9CRN9V3wSFWGA50U7NPweE4t8jXaK6ezMFFx3dL491fTgIal
kRDrnL5NIcD4t3HsOzVJPiw+peF7M5o6R9ay8XDEeikbEuDnJ6jGRPgFYODz6O91LO6lLaXTQ0ju
9438HPmsaDJD2005hTB1L7TREYdZlr9K6LLNx339OLF8E+SiuKsP5D/ZONWsK2RI+t7djvujFK0d
B2H2yqyoWgujZEqzCyQWPdcP+7togKsbGaWbuBzVKyIc46HQkahgS8zTTb4yO+NZEnFtbceB9QLM
Tqjw9ENGGVZI0sawCAjdLJNA9fH3Jn/yIfzNcrMGtTmX8P0J+rQ58hKSnCM+MCDG0K1sSRCvqpeO
u4VwX4tLN6W4u1C1UkE4SbLNsK7Scs6n++XgiZMjzGvAYd2oiYpcU2v2JF08Ow0qOMfC5GnZ8QaZ
1FFQMVLySaWptv0lQ40FbNoKf1FmtaM4WQmwisg2etNLRBc9MEHhyaatevqDk784YY8Aj33JG2MF
3hGEPiRLRzeubz63FqLXANyhK8ApKxZ3ywpP5E8R+i2cuSLVwZo5FFkljqiztv5dK/X+DbZt0dr7
27He7x7zFnrTi5ba+Z8iZIh4uWgBZYM78P1pKZAgDAwl6TVtZAWTgGOJ+gTNFafdsdeyswtgyV9m
fWzkop4doNS/PCXteLH2vkA0akVHLP2vq1bPQ9bAdxdnvSUP1AS2evQd+hsbrHFxvKXpn1ohtQmT
q3fEuPRYdxvMD/5LZSdR1m5nNbPuEycKH3DgJtLXQ9Y0p4AoQV34f09pdChjFMz3YjQvast7Zygv
jg5GruUfOisEQ7aK7eKHRkP/AnfNriGiUIFiIRfhY3Ax2KvJRhR2O51LEv68bMQos3WSSFQSFxeH
xTiznL1DWado9aOju6nLH+qMS8V0kfD/AJahG7iWf2UzlF8qzMGKe9YAEJw5TrMut40elsgq7d7H
QlHhkPW/IzhLm2yUgf3JmZtbyyN0emyjwKeHiV0ywVsHFg7Bo/zYBo0ldMigl3mhR4bYK5fNVsqJ
nx8gfBT/Q3/BmfzXnHMQNsCJm+IMva2YMiUAWA7/nWO3r63WXmMr03ZFXZIcjqG2vPpJfPtxVreJ
UXOWPpU+20bfvROwX1eiDFexG+36wx5JinqC6YZ0YXsBfQ+IzT14M+WBJ9JDeG6Z8mrh6lKPKx+P
HrqKWqi0CHf6DFvY3oCsvneyP2/ZBlgCAmQmRGngKbBVXXKkF7K1fC0AAaJOiFIhW1lapf5OVieP
neN7LgD1gi/wfAuLropLEFUcLdyRW9xyuUkFJMf/x7bcPJXarmtxoiLhRKZuTQyViax1iztkDTba
/2eNFD6aAT+7M8+HLjWYTqpKDJs5VNJ29VjZGN+u4ln1PaZtgpJ/DTlT0Cj8nqGPqcxfcST2OHMj
THhxSrhlMDLSEv8JF3jWkltN537XzeoHv7UEVSIeTyFgb9tPIS3WL6bThgCRsPExMfgj/FqDVosl
qMctLmIFWw+e3nOpTqHp7GQxaETIqpJTujB5yFuO3XxeqabekiyqxR//UQtScyoIr0JEeiaM/qCy
YUDMv2e89WSvv+TqF0+3OegNL6ENhkT14dyHqKihbRTe8iNfuxERwJLth7yb3b3W7triDF0mbZNJ
AIxbcVKCDQy7jCpTSIskYdzonpIH
`protect end_protected
