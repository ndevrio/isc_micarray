// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Sun Sep 22 20:49:28 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CjLvBbjekfZwCztzfjOsBvYKomCtAY/P1bSz6oSQiKIltK5V1YDNip2VH0pnmHVk
Y7+CtWPshjSbEbxExlN8GNEAdCff9Q9rxY9/70Mg9NGWB4vfCAqe50fMk9TT3PrC
Ds/mwHIXofB9avnVZFewUnEkIXDpJovu93mbaMZ8MkA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16784)
glf/V32Fv1tieaj08kDelR0LWAw6SEDNgG5B9pFl/KClNGSNlmumkFV6+Jwn4PUI
DU1dlxBo1V0juBJutGGgemQ5w6NnoWfbu+ltCDVFCEoSUNdiAeB+FMI/bEe0X7Lx
vJkkxX+NrarKhGPqthExZ8/ZK3KPEVnqpeh1SDBN1UOHToL+DJMZbFgfh9MUkOfF
6Yg3LMk3uZEMVB53OHOJHvWH5Os6J+zSPujK4MyeJvbu9+ibmaBpn4bXMpxC/4dt
SvamVNFCt+ka8sFXpSC5o/OGCTCxzZPsfjdXaoMBFzcnwCxMzKU5Vy02qNgB050I
7ZM+nici7A6m4k0wej5GcF9WgsUdK010zOvT8Yl9z2hEnwMi+fEn4xAYibgF44sS
w+IWcZk/zAuTTPrp2N9Is78BWzv0DjuFns6LNvgpSefbShNC/JW1DsG0z+Wd/TVc
C6dVfXsNfNXGFPq5ees1mOC6zYhV3wMVL5RwReqF2MzVyAMWf4Ub/Yk1rOrCtPnC
6APE7lyIwPN/plDSN3jPNVMsK0MjyeLW1tsK1tzDQCpZImAmSayMdldZ8C6SASK9
QpGszm01KEa+yLbPYLTVnf8HuJJvPl+cdsH9k6f1Xy8SnuIV7MGX33fSjpXtIeAg
PxL3+JVFcjll0Y37cH0TtFwMsakcB3G35W8N0vp/qnNVGJGEiaVjA1J14BGV8W/H
ZaeXTuDCbYVmwrLEqCFlXVD1SHSmAGPCec/TlvHKfbxfzO3pGqpKeJ8/FkaNhGQY
LHi8F4TEHW6MgkGCrHr0goK8zffp1FVxgIvOfLPii4+fd7Jv/5HTnaHeXnA9Tk8H
AOSnEWOaXx/SFUYoVyI+xcWSnUpRdGFjpzcYK2ovaBYU9OuNDRL0rUdwjkbcPgqI
Hywu051ZYu+c/RQakC5TrffDX1gkf0UFyEjYSghMYe3bRVu5uq7KSzsIOYfAmslQ
VIs5IsWXa4lcHKNuhm6FgmWDdc32WUOQuvQTUaNxDyvHsUh8up9MLRkTdaZUpObH
nyiaBGvir23K5iPT0qIiiuDMwroSgrgGoGtZQG6CfHbeRJhSUBqa+xFE3Z2ErLgD
52gEftgZznp6h0fVId7aSTHnKESTUdL+aMiJ1wrvOQKRvPv6Xzjvnk9GGG2XSTlS
1DAQ6DqwPI9ca2ivxmG9AE/nJBBAbUUcrYwfpEXLGI9x+2rX+HC+FwTrVDfQgzG2
4T04k+JpWL45d1TXfMEHAFRaGl2QZvOrYNmZPEviAuvdMWZvvlMMU5BJ9SwvxfVV
KqWWuDx4D6/xqxEC9KGdFWtia3txEvFMrU1Rc8eKQxUAGdZue05bYaSYtQ0hy7e5
DULMQ2Kc6Nm4APbmTNO0nNOtWFtcMIIpdjDC73LU36ws6Gkwm1KuST4JQCGBEMRV
Grc/MIP48KqUlh1lT+P2jwPlGnv/2fiI/yaH7eXdmPUtVoBkU2JsHc3au8o48QuT
zRejjGG6HU5eoUNCncj6SjilZtelCs1B66WOVLZg3mYtCxMXl43YJ480KHXAOjag
oG1F0mLFtyhfganMyH9rOkP8RsUEDZ1sk2hJJpidJ5qu2+wEtuY7iN4lF2wpjloh
7H5UDUd+TzQ8tqJUaqx6nz12Avt2hnvkQ6vSCtj4MZPGa4KzMvuv3ttbVuHmVbaH
FANzb3zkTo6Wtyu9f54GOOb5PylZdJpDWIAXnV03B1yhlIgBmzJGcHOnTsp79WAl
brMDO52QIhg6FPYQ4EjeVlavfOaafdJGKrzc3VpPAKi0IX/jJ6OvgUS2n+4siTQu
NE5vv0rcyCNdLGwvc2BXEbUGtryCqkjzdu8Lsse4rk8hqOl388IKQeiRg+V2UtM4
PFyUH/3zIQAbR245rjUSF75ZpDfCQax5haOhDFNJwxy6cuLmnMs6OMWxgXgr7+Lt
mopahKjbHKKykAyVLFGJmHKHswXGR9OaNNie1/5iKAWRp7ulUhweF5amxc3+lQzh
rL8tMG/g3SwRb6LT778NExfzUl56qTYAHfKt8gj/Ph1uzA+v8B+FVSnNfMPLnOZK
xL17Vok0EDvDK8rSYb1cHmLJEeVMiSX5CXt1ixx2pleL2K5GNCgionUTAIiJUNo5
86msmwDKfilJhWaBNobjp8L9lUwHJn4Vk2tt4BG6A2N9vZ1KNkOmyNFrjUjQl2rC
IAjCm2xA1tFmqnzipPSPDwlcMkbETRgva1nYo3WY5vyoHDaufBxq6OyiYQRYyEnS
xzKZyHYNlg7GKDRum/7TfYLDO4qTtEDPFNinU/nVNgA6ufmFsa1qDR5XnTMNzUZ6
VqtTZqj7HjcaeM04+OOjVneWfvfBNHFop13wRUIVSu8mJhhd8kKLi5qA9Z6zcZj6
3KSgqJI+iGA2rjwv0NksKjeQteYJS8coON0Ftv9hmsntbb6aKANcjuQKTNNtbQxy
yi253l+jsegiqjJM9foDiCO/zzb+1lTO8gu9zUvkatR883RmbclXL5B1ytzzXM8L
IIjpjDF+G0GZMsDWyGD/Vs1nyUrC8L0rBjTIEXRlAkiHvXQsT4xq5TsEA0/MqBsw
S4LnR/e7So0tx50xhR4iBmn87QWc/IS3XDyoSsXfAEEaw+rF8BUEZUjMDM7Xgstl
b2NI5K+wKB94rH0lkEQXJjtPQfWfbkjiywDyXPEpK0UAwVXYvrka4xMh5rdz+eMj
xpyd61QOZsjARRrAs4bM8dFvrbjCbLbhXGuMPVNv2uzJE51gQgOYlEy6WCh4/CkQ
NXYdJJvoQylKmRRgSMw4ZLMRhWrxjhvlWtPu3kxHYzqMTy+RZ6cp9tSQ63mnbs02
+Be2lnlF9oCMSysRN2GiKgTyrGYmweNtZ9zTF9p16+SHOYx8PwaGOUqz56SI3z5U
OJrFalsu8tmBxa/umocPoTTD18NYP2OzUn3ZpRc3Jy7TocGB6JNMwmEGr5xrrgc9
Z84UI9N1PaCVER7JkHVNWxlSCgdf41p+q+5gvY7fK9rUvQiOHnq+bffCkBPAI1Ut
SeV0yNs2mdpohZ0lHUo3pWUCZs94mABGJVysmnJQ6EIRRd0Ee+AfjZYgUZKq7s/n
792jvF9tbqqTvcbI1xEeDDZ6HZkGkxzPp1YGC5buY8gxCxry66KtFO8FaiY35x2H
Yq+duTDh3QrMBjNnFQT3cZdv6hwShI7F03AM6Yyp4a7Dcd0ZA4Rnv4P1OL++ZHyo
TcU02cWCr/5vzuof3k+liKDMeGxKjyqTr/3mO2QOsVPpxwelkr87XmARdUlqcydq
9fOm5Fl5BKpwap9ZMK4TwPfho4oc2Zg4JD8gMO+78+h/kZnxJecsOPxJIOnkA9AH
3YcJu+j5+qMAbW/ka8RwCqLAdJgORJ5gZr35wAzSWYTPOmVqiUP/Irsnow5s0V8p
rg9dIIOMS6Q2k+PyZGd9XY7LEC2HnBxTmZGd9yR1fDVHnIZKM9t5HEax0QVWvexl
0+bkhvkCR6W0Z9RiJ+oNqpU275SsJl94otioEDI8K7lkpOc4HuaDq1Slh7aQhaYU
Wc7RsfUI1ERCb+7dgpSz3FK/lL93qazv7ETOl/TXM9Lj5d2DDWVqxHYJfqwqT39V
RLPL78xpAxp4y94HzL6QmpY7acJ9BI+1Po3LlNEs0YQ/pEIfeKFJAsyYTPSLsi8i
i/tcUuc4G4ee5nc0lZ8hQfezo2OrhHZWsxk05iE227TSgr4QahFIoQUxYTYzbfe3
H3rz1S7VyIfPnbRHVKS/s8DwBgsFPBUSTtMflF2+UM2AtlkWoZ4xwfxSkKis3jTm
5BEvwOqgEbS29AcJ60jNUAK1MfDnYa89inBMdpBCHDCnA8+/R4das4rhrv8Ao4VP
RS8wQtW/r1aPMKY0m1fLhjna79wOq6fb0rrQQsbY3R1WC0utl5jbANWD7Ax26JMq
wd+0zfbJYRmMzEZ27J1NvhoMjrTf6/3QCArgvcXOfYkmuQhvCtikgj1Jpkk6q9s+
USciv1ctMqLELhVJEhOnk1S/tBHjBPk0bdLjQGfMFxtz3Xiy7VDdaYB6VglEWJgY
LjcitKTt6cYusR3PQ4noqJXKwP/h8Em94LhRVGTJT78P7gDq45MILGADtdrubyLS
NOsVPPmIfSMcrkDgQsPck3oLNyksRemfHsWZz3aa4a2aQhKXdD1SCMll3dSUB/v+
/NZHZIG573nix4tH5I3e9fTVlHQboAG23znF4Xrq5RYq+9kBMAD1B0G3WCJxwp2J
9ZcgFYqtofmZMc/schtUZ7GYU8vOFN4gGnXz4IyJz+x4cTKhrxXDRBPUZpr7oY+S
IjY5/OyAUAcu1DcET+f+Yg15kZRXDh7OeVdcLqqJfhQWYr5WBAp/Xumy/nTlRCZg
rQBDZyw2AdiP7r9rIPQ5SukW8zKImRgMBLhZFCLJ+6EIIVq6rUjXkIwfiNiwb272
7EbWzXGUhQp5pJio9I9CjwxF4XoF/xrTLQzMVGGJsnFJjZyaoI7KNofz60iakMlN
zBNNBqejcjlMictj6kTEcoEc4h485UxQxz0G5uWFKSl6QgvKoCt693p2eGEAzKWo
zQ0L+WVvpnUuDCNX5fy6PZoB9A7Hh2arOlpLe709+bzk1oH+deez90ZsVDulkleF
90QxFXi531PxPDjygkIMbBFlmAb7TKFO6TvWY6kZ4jPxZjB4n823rpHmVj6Z787d
MxPIFzteANVkyqBL70TR57elTxRvskRktDNlr9jsIIdOsDqiBDUQpXmJ45nJ0cyr
f1XPkBqUwERj3uHWTSl93flS0tjyW5LUVma8ClFim3ii3PqbmqzHZJR+7hQYFSg5
/KBUOvWibobInQagmDIlvd3+IiHLnJjkFdoxhX3hyYyNg8qcUP5z6zgHQDnKAm6U
cDR5yLD+27hPkFjyZVPteN635yQ5J/LjdK6bLKoh26zZD3FW5K/UeuZtQM5YsEQB
Flbmb8bvMF3wwKg14/FOjrzT8O9E/D6GgItLcmGvzW1OBVdQBV/TybVqZPnRrcXz
uLgS7fvlw1zlBiXNQHv79GWBryI5JfUGVMq0ne/zaIXxsEFMSmq94vo3Okw05Lsd
ZqnalMsm4xFLxsxrIn8oIIHnuUFIZtcx1/j1dU2OMVgGPGMFXhyhWkD08EzcUTuF
EeaE6x3KHEj5XwYdeK1CkC81C1nzcY5ReiDZxzgMVTFmWJnhUtG/h/QnQRs/g7lu
R9KK/GJ7JyXIJ8u6bxoV1prMbxvfYzESSOY7i88F6uJM67+mz5rf7Q7lHDL6ThcJ
w4uHHZbdwOC3X1yvd+ISrrimiiN23aNlcV2PaFOtRo0rOeN5qawYYvAMiAth4Y0W
v+X/w79shPnN7lChW4sdzGMfFSbhIkt9sfcdmQNqpjRUCh7/FUDcQrN1GjvYSCvk
8/oIY0FCoaK0ozAGM0YMMdG8LXtguBh6BXIY+PdVvV2+W9aAX7RyOynHNGbQf+v+
GHa00Wv2b1Y0Vphtku1qjcRc9vQturOSvkB9cUmBLRUXE857GdSEx2XoO0wOFcRt
mclTSwfWBL0nWVe1VYtZm5FXEcKPDQGRseTzbWyzR0AO9PlnV0MfrBt865Pcemgq
gRfArIyPKfmZtUud/vt1jZMdsicJbbLhEylyABVEXwoPMQNCHZ/g9hgQQhixVm+L
tOQfKMdcKBo1nzrJsfad8OB0TlZrlwyMsnM3MqfpseMRmrfYZxtKG8p7R4zBDGvw
IqY4BHXfhHsP23eQoUHMiFrNklBtqByE/kahph9mPC2UlP0mQcCO0OWLlL+UYknf
IUBv//aaHPdu5BrusMCRuJcNv/YaWFXLXjVeBaxccSU0zVm75YvDlh0wyKfClKd3
hcXh+CeQRkJeEiKYszJlKHqxjE7Z4BgZ+4q2gckttsZD9LHO1wUzveC31pmXcldO
xALYswsJ2nin4dPjxYYFvQqkUGdXJuwKoCJ+u8JT4SP8i/0CJ09j9Kjb9GIycMp/
Fpe9ouaiK7fEgymzPoGo2LNqKJ9ff0UrTkW4jxGwg+oVmUwj1rFbWlDeTNtqqj5y
n3zj9Va2KveQ4qRFaxaOBHbW2dI5P+Evs8mf8Kz2pmyMxVesHUi77MedKD4lauJb
bj0QWSe69XJBmV2U8+DcBfy7Zes2SsNTScW0KMLFzg1GS+A0rUQMNXmDalus7F0k
PuSi293OEgxaE2OtT9vab1q/ZMTgMMTTJ0FX0qm+4GYI9zfnMrOIO1PARti+WmCK
91a1Kf1I7QFyRBbkwlP9k2gdGRnhLaDcUUXXh9QEah5vsPFQfL7+kclQ73o2q80j
76UeUoL+AMuWWXv76wUJLESrnujVBzSqwXDFGDpTG2z3EwEQY3goc54WKoqhGtww
TrBfQneEqyLkjaLgMRRmys8Gh2fWTkvKCulvSmI3V6IDTUOmv1wkjrVcDdPCvqn5
3JLw9PUxKQOOZrte2CcDqdsApIaabm9Ny1YEiQryWUBANxyagzJWGbl5BieGFvZs
8/9dRah+eiikwEWBMcrD55tujnMkg8dLi3jIAxnXBMd87/upa7BfVtcC43z6aU2G
3rO1UkAGXyt+jlDnI5vUS8Olfye8ihZTIQUzn8ZwHWiQAr0+SiiZAYWW0zH22A4q
sTV6WwETGAG+Pc/W2RWNDiZUNg4uuaw6YH6DlsU/lRJkqx6YAOKBPeeGTPMeq9NA
S2i6BZ/p2j8AZvogbAREUZtsNM2I6u/X57gw5+xIq67i3KdeZqeRz7kvyK9iEcpj
rDc/DI4C7Eqz897X5Kjs6IPWs2vDz3XSaNPNA2A12jVaYp5QhTKUKYXpQFvY/lXk
XQbxcryx3Oc+GKQ61yOuXiC2+2mYjUFqvW+FEY2DNaeIpM0vVrBMC7uLNZ3Jcm7j
70ymoxsbGzdjL+tZ0xLsIl1cuZnxBLSFQc7nGdv2P/ueoGbtzuEp3GpA9nVwpBZd
sLr7MrIBQB7bPo5uGm9P17SJZAQNsYsSaDN4VwVtR9u17i5Oldg6xQ+tuOpDQfCU
YqA1JbpdHwXMtYR31bbfaMliNIzn32JJHC+puZvomZYpXJjkPEPkrSekem1euMx6
wnZVwoaiZa8NIFj5lXPCKk66OS2oepMM9HSd3Dp66359Njk5D23N2a01DgfnazYZ
NKpOqODhcah1KuxGulFt6l4mF4zd+gd3JQK4b5QzVt1FwaMD4uHukfLuP4ZZTJc0
cTyGJcVvxbCIVIY/9KT/prvu7wPPAS4MN9JpuC4/GqsEcnhv/HMpZLnKv4SBN5hf
2vIVAWHYXvl5mKjcMcSYuvMyv01obZE6jwp8YZ6ri9dfuGYIEPkxK2WrCHrv3X+G
yTD3LEk4c98kQr4fFrQSIfH0Dqv6MELUqzkMZe8g+YWSogyqBx16RwD8ZHA15LJA
MFaX9uUIiJOPvXUw3Xyv9Z5Ghv/i7XStMZXXz3LdMkLgoUD5dw0WHT1iZG/LSZoR
2KbYWlvRPasNCYfUi+o8SaZr2QBVEPz8zn5YI2gxm2gEFbYVO9jTNP+Pf2lmhFEB
UI1dn/EszwbTkX8pLZ8FNqEiVYEfu8xZV/2oiRDb2388f+3ZybDe7zCWLBbnZxYU
IEK5OSipVEMzWhou7X/VDcLs0F+uQYHbFbQebvHNzMBXIlOGvczlGP5aFS8LqaJG
m2zQr9WwGM/YBWzT5jBxTuT+jgHPAKwOXt/SyUPp3IC9WAI4brMgV9cKl+snHXNp
zzUlNLzqum2RENJYns6v4eYBW7ezh0Eh+5NiURNInpSTyFmISceAlT9gUR0dqUnh
ElSs5dBnAk5FcR069JJ7FzySMLhsEL+DuDBaUyK8j7CakvuWct9Jv8LpL7IjJVRE
MIKi8fmt3tqy1ZouLIGQ/b4HlVb1aS5BoofBs6RmxpPwELs+FRRqHQ9f7Enty9lN
OBmLYugWprFY+7dJdZqRXY86BM24ObnspbH6GlD9Vdlm/CBUxOk5DMqSCrV7Kud+
OvZ3YLXwcbIsL4zljcoQu3J8J9YpAEBGOQEIt644c0jI/hxq5UQM9DspfSghPYhG
MIMIjFwF2/qtvEG00CmEjMexM3qHiG1TDcIpGJzzYnAt8WTBMvfxPdyfqBMtMv74
771oFtLzECLTfPumIJpA/YBDd+0Rs/P7ap3bZ7HnXy+HHkOhs0+ZAxnFIovN/qXL
1PhSggPnBU9+i4bf9Ex7PSd4pu13WbEn4KdHw8f59KaKpSntAJHI+ngXc8c72dT9
Z/vYvLm1gECzapYKHFPODWMYbJt125ciZ1gwIo1NC9O03mkm+7z9doPiee3+A0ge
gRs+Om/SvZHpptnAybDuSPWA4snuwBiarqHLvD/NVEWiUgxAIi1QWe7bH1Rrxm5Q
BUaBWQ99GwRqvrqEjyFyHistzpllqqfR855aaFeS3K5m3+1ydppPTpmFOVtDw5HZ
6L1prdvAn4Fi35GqPZtXYLoMv9IYtPcR7hNQPpb+uL8z+zTGbU4Q3NCPGNdxwY9p
O+XLm5AQaYE5j/CPC4VD+f0ejFw130LC7I4inlgqbTesKWnUYqxICZBLhZWlXWiR
8/8Yt2gI4qlQmFS1+DMi+LtjjfkzuW0NCo5W+R8+6u6U21PJAbUsjScpl3ACkrr9
kcZmoHBCD/2m5iQy+qSRj+DcpTi+kpWUhiV8tA4Dq5xhTCJ3UJc4QUnW+JgrKWQl
rwJLLJbBAW+3V/3I2O3tHJM1C9zCOjPR53ZfNSc/aaGO3eyjxxM3qYAQdIe/j0hS
ot/WXpUaIJJ++NEH9OsdTrrkdVhEixoiKU6g+Qgw2pFMoH61cWH5pZLFbNd9UjSh
kWpB2RrHSZLAJ/9VcAjfyFyDUg6OI7Kr7YI6avrGIcSiEzxfsrKstjV7ekQcPHRf
4ruccClCeE8sgMLwWmWytVKqqDfyRU+WkS2PoOLkZ7PZURVt1UO7DgnRZWZXNB1+
TV8rY6cNivs8u+mM8fuiMY49GPxQbo0TEG8YIR4zpxYsXb0DfoUMdYjT8a7SHixj
lKDu/AjNy8CIEFJiibULQ5JM6WVsUu6fMtdOwlQJCFcKw04FoY0hm9EN6kFQf++B
b8x8Va3Of3ZTP4QE6C+JmrgeaJdV6A60Bhox64/U/EiwN7aCVIBalULtW778zu4H
TBOW5qa8VqZbOpXBFOHNY0SLhmodQK+M2y3A4G0rZVJbRB4P72lj35F5EaskkdhV
CMVyP3xvZGxpGAN9H0kHmswp9s9T9a+TeEaEDzrHjXBjPkts2v02Q+VlF+JfMFmt
Pfc3l6l0VfwKIj9ncqLFwkPKMcZbB7M2zlUEDzT7z8doLf7MWcT04f1o8S5SPAyZ
DbjkniWwVXxraWzpdFO24j0YONYUG1aWgVnpjaWNUWNoFoGy8eofsA21HNAqfpFM
fTLbF1ezuk5R0vSOHrO0cQ/JspviRpg5+qumveqCHXj95/QBeRJN5YhFYNWahue0
vvfSPrxp1oR9ojRXjapw4HAksVyJKJXIXbpVnQVzJzPhhE1Hwf1iOnQdn4Qadrfh
TBNep1AP5aIXs9myhbrlma5kNSROmfb4HSCIqNjTPrFuEEj5jmd2QA499sU2nWKM
Cphh1HBDzQb9p0M/xtOP6/mMW7TOb7zU+I2gHD3uPQnLxsa/GI7Y0Dg4eydft0Dg
U4H4y+YRxmTtrruPoHZY3ytoM8xutjtCiFrgW0qe1sz8E0qWSK0j8T9rJKpq04EL
TYShyQRZ/CqZViqrztWgBiQ5XGa+lesvATHMLPDJDghQLj08UE+d5kaiSlxmxf84
+ruTKoHZn2qULdimovKybr1GtKbAWxjlDQzqAkqFQeSC42MAv2ErDPymeUOCZyMg
amvkPf2eGSrcBSP8jX3tCYfNlq8snxCICW/PQs4XL6KTGKY6H+XufMloOQgga3HC
S0X7Rq2MakMkFw9Y2gusPMG+6SG8KsO4hgnGE5qNkznrJxY0L1RyHpEj5eog/dbw
pyX5jFmkgbBAeEY1pa9eGzwFwz2iTVWJ2cR7Nqp6U9zc4K/8qyGa9LnMS4pPqxv8
m6ufdS9X2lH/qG5kdh5zkVXNzZl0V//oFHnZrWRALRy1PAhXONZEHudd9s+vnvD9
Z3GPBrTaL/ArxpSnJhEBile170DF61x9e6di96gawbLfMdytHc2jxn8bvRcT5JTl
MkfNfJvIOqVxGf+SzP4A8Lu7IcHTMou/WtqMuC1RTT+5OcMxzBAYOnkTqpz7kYse
GaLAN8KZVvpdzupADIv4waxpdaZ7WVN227o8YyjyT0S3p5rfGPASBwoK0S2LUG/2
Dx/XRzzKWeO2ylJjSUCCr2EQbNSYQc/ynBJD9sSdHHCRiMRO/prST9p3wLyzqkoi
hc7wyX3jcB3j2y4jusO6/Tw9P/UOPwm9GJaOLg53tMwmNvyN7pnKn6U27K5yOjo5
N0Hk2aVZNCo5py9gxRnlxb6ZJKea3dI0GEIexGmCvFPySx+dwvCmWRN08OBzDI3m
dCVnQD5EbZuc6kXXyM5bV7a4A44sbGPjjMdJ6F+LHV4JS1uAyhqCOaFy1ZccOYTb
xTeihrkF3bQVnAxzBh5QxnORszs7/6B/Ul8N4fPa1/VHpyQVWcVd/I0dmzpP0vO8
TbUBG/3JPoEaDq4RpQ2eezUH6Ln8NMIEhHOCrQRyUTDWF6Ht6y1SXXMVJIJ8+TRh
Twtxhu2nSRVgC9Q1UvLDJSIR1VNNR64UismOSf0xLuSbGbRXFJWWnzxSNS6A/Z6S
xCZTLAZD1kN0b6Rkz/+/6KJ3Bq+IWx1WIWzEJezndZ+GzqffPDf6XXN+OH9TalM3
GDkdIDh4ojhf6v5dO/NxtZiBnGtlu+BeJSBxpYkAlPXQyIkaIhCaKJiPYZina9x8
ScK3RWEkl75PId4ZM4g4bBMaf7saFQoE61OjRqHYy7bROo+io8akzKkGsY2qqYTh
F89Oy3CJVBdVT79gzyY4C63cBPAgQiIUFQDbyf8Yx2I4jMUQXcAwXF9NNe8LgSOJ
Ccz+Gp7CuVK1PbNXUks10fsn6yNmLkQO7pXxPLc+oIncuoE2H1JDKRvI8BMDsLfH
bPuRbQ2BkNGXQCz90Ur6k18/UPpVK/D1sMgM57XOszHgLWnD4jgN3PRuDs3VFqed
sHqTVG7W6qsg8aSB5Cltr0q3FqLNEy4bt8fQqVTAL5ctxA6GazytCROyh1BKmgOV
bqn6N3AXm3YIXt2Fid1b6NLrw1wsRggB1kxs8zOAMSsNNBSpsZ7GNr/P+XoBboL4
aNVN10Ru0aOOhlDC/XPxJ/99/6wt4JfGyr5AoPy2YzJyPrV+sRQ1o1k/KoL6UU7L
xjUGYKepj/7bSCG5PZsPn0tLc8BGQMApSr74IC0XSddSNfNERkxPHff+hlqCj6fo
el9Il1635VyaMQFHy0Hzg37hAHXnYxr1hK/oiIG/0p6JqQEV/U1xHfnw0jSPZv3/
+egELaL/Uk/nwkSZ3nONxg/pQhmrWCnQsbVS3wfamDPy1JXKrUT4pEUYq1O9fNgo
EfPwDn/n5P2X74KpKmyrSYp80Zc5tmiggXR2aG9PeFtCeA5OAMnnzaK+tSW97pEU
OLRvIemBl4nGNQWCkA2jXGfD/gTv4tU2biBhe46/3Cd5bAi20S+J8ev+jWI7bx55
mmPeifM8GiyUFQKZfST72Zeg1A25niMLvbVX2RwLgS743K/FIDRAxG0BmfOqTzuL
QEmnY9Ku3K72dQi4Gj1/pTs8FesBfRy63B35AE5fm0HuYfEs8Qd5ZY/J71pxnqYw
7/MPRT4DQmL7HxmiPonPzMj/h2O7/XlBTtmhKpr/aCbYEmp6Ox/DodBNRnBANGDG
R3+G3ltcZOotwI93pVhYjvOghNgp7uGZ+hLoYcd0hKldzwdYsh2c3P3fzRaLENYY
ci89f4OqnH3FZucXMp7qub3ZA6cKJE8MhE38Vj/UqNqqyMptkmV1bl7mVufXjWsk
+lXU7DBMuxxzN7uVmObmDehhUZix9rDNSODO+Jp9TX8lj9sEAzBEWe3R2KaFYreC
P2H2t5unvN2rSvF00MShM+VmROnJWivkMbLYLugbuOzN15g8WbqrAFTfGK2qgpRd
n43pufYZ42YuXfDV5b/hF7bJiIqNxnrMgkFlMPXtzYjIYj5ZrnwHOp3lDmGo+eco
ZW5whHr53RZhkf+TQFiu053OCtCrkQe90p38AzWwGMRgjUxJ9pzQ6Qat1clYA0W+
O3jsETVoHaR/enXhJvePeB1gvcWblXlT7x981xztngo3N9Eiq/ARNVnwAp6RU4w6
QeFwAxFRVPQ4O6OXzqfZrl9RRRwM4wmVrVBCF2SK3AZJ/Xvp+pn9UfNYv6f992Fd
eqxE0zrgqMbvnaPo3EBU621yswXU28szUvGyMB+m6o66zL1hWl44ILFnS+lMqC7q
1/FFM534xAkinC1QJhEXk9sFfbqIlYUiGiN8TDYEnqb75jeHO61w+Qi95sH4OHJT
MIZXd+mVRsnhbQbA+wxVrH5wC5x4pbvMMBg1JuPXdphJVofVQEqxrNVgA6LVNvUt
/xWflNKwlkXPNle4+ApbthpiAiPMlUKnlzTHqqS+FIJE6ULyh0X6cyQcD+vZMLKf
0ha24Pv1YcfMHyWX8AAFSLbNqKHqKzjorAJmciUPzCvFYymgAf2uBjQCcHFFyMgi
VpWpv1sSmSQbRJt/2Xh8PnGooqhz/rdCo9jPJu7x6jKKBqyr9wRUbpREZ5a3NrpL
6KODALZreOQCKdif2vym5EwzUy+575qzLY/ODblGgeSUbj/tHqJV3Lj9ICOZCiHe
CX8xQ2ahe3j5cS/ZIMOZW4cruAoqKFve4zlIJ0ZPaHVpSMbo+BYONKvJ11CDUxKl
PP+9CtzRw4oUlXooBFgGAkfn0y08hCYpzcSVno39qIqciV09JuLvZz9MR42zlMzf
yir+qljHSK8apewqIORycMa6oE9oFzCmG/EmI4mYoGfP+LYh+wu2BTEJLNe0TQSi
izMNtKK57miWhM1zv7UF/iJ2fIPluZDgbrZB2L7rNl22Y3PFrG9Y4Pohzmm8wuGJ
oKwDlOYm85dXwQeJG3uWOJ92wV0hzphiI97BiRo6LomW/a0pt9gd60ElqC3vkh/9
5KqvBNJ5AuC4RGLSLLskUZY4wPyw+fnWck61g/AMnr8w3+wAhWjLZyeye3eLPj/r
HwBdoJCElaMR/U5vsfD3qBgXMkYYFYxNodSFWn4M0VQfotbRbq8aMTDB7MeoyDZz
FpKKeqZiiNP03Ur664QMyOjVqHpTePli3NdVh1pVQ6GqX9Tq3Of+p2kmKaAxxbcA
fPol7tbvgbUtzENJwQMid93vKvigh73XEkeym9BCefm3M3zAApJQkcWtuxJZaa3T
HcoqT1PKUrwv/mKXgdJy7vm0bK5KIleRDsd2hnVtnmX83ixkcCRElervAZ0bWV8N
DwKvav5jWkGVGfOhVlpc/LkZPMmx/dK5Xmax6jSbMJ+e1ewfUsyXicQ2914kQei6
3BEDmA6xJG1CRGRHM5Cow/TcigLBjnkq89DcX3vb9GY+i3ZlHWXGnBWqaSQkNxq/
ndeUfuVSSvsxuSKtNFWz9CUr5xFpzDQFf6upriPnWJ1s0keZtYs+W2vywugL66v1
dx2Huhu2R/ztr0NAf8ieyEqEM8VyBJOxFFtBU9wm4TeOnihbxZBcykggoNPhcb1/
KRln2pWzDCnB9wUe4XpL3OugAkivQdDRVfH3Miq7dL2zOLxHsXoFWU1ADtAyf6I/
6Usp27Gc2WHIHhBOAPzHK5eLX8pZvM+ZG6yvSse45OFGz6NtSkn6k5o51y+t5lba
iKGOFYwILlgaQSzyKYt8y7tb1lb4JjxnX4W9vlZWLEXldUwG8vL6id0w/kdQhpqU
GJ4SDac3jtOqgP6jDl/MQU2DIkrbsvmTU0gTa+2Vrpiz1Fnm2ohOwT/BPzvxPzLm
Ev99/W50MGCYMxjzDK0h5i74IoDuL2qiAxYOepzZ+eLPCZ3Z4omLwotOfjLdQDYP
kQsqNS/HWMknTLU3pg4KVjGzTE2EPqT0ynRN53u4zEgiSdznGlcK+3qIoB9kOgTU
pYQGlWOHEncbHPovFdG0Q4fvMJcn6h/sPF+tjYNXjKL35Ucu9fT50GLuzkCZ3HIU
m4BIuJnaFf/HIJ3L3YzVNJkRIQgcx6YrKeC5A8112heDSruNjSFaqSAMLRiHfcA2
sT5eKInyZs74/j78OB7tx1a90avvpd6/7fZ/7UlBlSsG5Zq4md8iGFG9SJan2e2i
3z9+r58jKIA7rv/vOoNGCYJrmpNUr2q2luyHWcX0jEwcnLCCfiXQlmmjilKqG+A8
YJNK0uGek6YTR9O6yRNuVHsXdaBBNhfK4uaVYeRJrb/PI3Ke+rPlM7Umcc255HVx
zBXUpzCLCC2M450Xx6h7dOptD0Sv5KfbUTuMYh1hFFfdLX1Njm+SHCEnOAA4I4Pe
2Kgmjf1llbeZV/T0TUlxcPAbeGlFQXdXNYwXB7xCCcG4fcrXQKRKyvzY69gACxuA
QILfLHylfaiUWcqy55U8l6Mjhr0b35BNpxd0c7s5JAq/EH9MvRgZuzjVwEfcTMoh
F1/sismTNb9pMS+iRtgoIHX5x4NItN3sHqzr4CrcjvXE6rIHcoBM97pmKvMmPHvW
iovu6FEe4+H1nMGGkpgpixgk8IdQrF9V1qsVIGZbUj+Eg03fat1JUBAZALW8ROig
TlHT0/HCVhOW5EiNAwAu+rBxBcZ1ZPvKC98R8DXgYMALUgPxSy1w35D6yrfARkxM
NHg89Pd1oR9rfOZVGtdH3AJ6Lm8vWF6hYwoPqEw72mrbi2K3SWA8cLO4AO+Kundf
4Ly6gfpr9dSex8vmyGok4oyB/RcKy4kxf0EgS5GgtXKRnXABWIfreKzNv7XP57/H
OhPeykWJ+8i6MueVlSiqP7RXoS3Uvyz0IAbnVf/m69toxYGjnJj04sL56OHTZXIE
VTaNEXMIl+v/GT/p6NqdqTbSDejaEopcxjvv7gu45gNqRYnkbvyvOjK8a1rkDTVB
Jn0hCwO+s46x/wcM2f15A5mKXb+QSduKXb0U6RD0zYxYZb/0twleHi7Z3iSObAoV
HlUxu6OKtyRyS2yNZfTF7cHSJkk+eoKfccidOiNo0PQ+bZkB6gMWdwUJ20YSwrC4
xIMwb1Ellp3rCZTpWaDhiK2RfMcGgnY/uujqzrg1zME3j0yljhoGDUmkvzwnXHfP
K/WqGcWhUGOJuKMAjU6RyzqRRoFeAla5LlkEqKEFQ6m/vPEHi4fDAqJ20dJCoJpD
GUQBRXLhbquT0JC1S+h/whlcXYDRzaW160l/MLWnsB7S8CKHCEySRLpClIFgWURD
WQHvDpKg6umCGIIhCFW6igL5Od28V6zMLVxXwwyvkaruSsecDG0uxJUujzcHmV3X
b5UE6XLcjNnHCP11MotYzl/8N0VLSmP3h4SDGIBHwKX8rFYm0vCOln7sP5aIN0jo
u6UjHWKPOtRNsKdtx55FhLQbPQ/jd5NYP3gki60Xn26WQEH/WAPxwu1AV9tGE5T6
lZw4wdTU2gZPe0YmzZ+Qa3sIiobTdz3FbSAugvRGq2nVbFewaHPn2W6w7rGtrbYg
X1wtKKiElNDfyI/wG4GMudHQOa8MrrE62WV+Opat2AiaFQ6DqZcN9bZFbb6gXgda
g/+J9Y9KZnkHj2UAvNec6XAHvq1YNaB7rvGZ5VPhgdrzpduUvlPCg40D1l88mqzP
zLF/Jc4asbRo5b98MD3Dlz4LCBhRsm5gX9/j5zyMVBw4Boz4doRkiSpn1YzU6ktj
6mTvJ5H5xVpqrU6BSefiP4y+eKP/vd4NcszDcSiR1juqvGgRVwx+IBEQRO0tbD7s
MiccZnNu4wSdxO5pFbnwTM6qz6JLWZGAUjmpj7ZK2Rl+/At7LSONECjSycwh19Ni
ZKGR5JoiSrBkQ/ne563IiMWKYp1fAXtUCpka1ZXlybrtL+eaj0PejM2enB5fYrqk
HhaOHatLzyHZh2hln0x1LWRb0OA0v1G+xRgeG/TmGErI8ftZt0iM62CTvigHGg0t
/FOGVu5CXpsxTMgstytcvKcD3JCDRQlxgd6cHtCUGXQYIHV1Wb5rmqldZ1nSKGnE
u/pSgD1WSfRCLwDZS+TGN5tR6YyVgowf1b/HNVcQt0g27XUdSI1CSjB9F+5Y3d0W
FdVuhJd92MS21M8pwsZFWQWwOiqnCOR4jnY7ZGzOkzgIJgOSlgyIsivy0i7YkRDG
iz8D5rCIIeYoHhg4iOAlHnoFJOitzPH5fmIpkmSTd4MbO/I2hk6ZzfXmBGUCJy7e
wGjoXTRpDtu/R81c0q+qCVMRpXzaDRb1+Y5TPwQaQQ0Kfc6GXLF/1Na23UBXxg//
eOM3d5DQ3DZ3Kf5nGxjIMSNWC+P8O6M6UkPsF1wS5+wcCK8ybxKjU8B27DV1awkK
D1yKoXbpYSELQAYXmF1J8glwLcBApz6yw2LtiIoVwo3JNYTa6kJQMuMBGZG40XK6
jDZki+cSLc7Jufd+W9tT7YumbVc9eRy01cxLkMzSMkfMrJxWvx9kGMdqtq8m1aHC
0zn5/Qvwo7TYLU3m3atEWQbAZ+GdKdEoryOq/XljpC7apTzNw9buRCw1xOuhb8mW
9zWlxYi9tq3VYtqcBnTJLXB3op1K6LzRZ+wiurJjeVNS8LvRrJgIw/lw8t8yhH/B
8oAcrAZKWczsW5UDPzKfr7eWVeT90KQ0UiHSGtJvwFBjKktroe8pelwkTKM8stHh
qhHOwznbh08qWpY5w/TGP12K6bjf0ZOrLl0nOf8rV5nukSbWXUdwk6/PUxPvg/FV
d3ooCdj9OJRDLMMHvjqXQrO+LiyHD+h1Z1i87UDaYmj7hg1BHHuWabscNgXQ9Zyd
aUv6HKmGO6DXVt70xlvmH27P5HkmYxJUOu7XClfuxJOfGgxyjYbmWt4AffeISAxl
eup6nS8Th/foCF4t8SD1TB/i/BKW4IbDEVoUfnVCYI6i1uexYr3G+RihcaCEPv05
VjVmV35IWC6d//TjpZ0wPtmQ7qQgSWd5OcjhYcKpBVoUxd5RyI2FHbiOEeS9OKnk
oQBQS2r1hjucQjAfmjjs9KjmEOsNHivMdc0zBZAubpe+vIiVTkkSicm+iAnKAflv
rzcgDdX6mzpfcQ0b47e8DvDl4o/Xj2sWmxiI/SQqvaEAmSpRYLvNWP/KhbAeZzh6
rkc6yPF6dn9EB0ziK5rLK/fG4O4NHHb70tWVO+Fz/E8oGt9twvjpEPe6XwLJAAx/
SDlDy68qu91I4MhzsTrjshGcOUvNRf3RkihQTh/0EQdk66rArC4b5m/D4ZWhBy3g
AaniH2fYBw++smiu1BWtnF7T4tY52vdbD8SsSYcdZEw8URk9ZRcxBrGJxRXMpkZG
ejoDNZ8zI+JzJ09laRV87Gq9+cn0E64yFXOawcufSgNm3qScXJ9Qjy7IH9cC1pIY
yrcFPqzTXYPEyG6BVpqpt46yOJo/EJT7/omoYWQ7ytHdqyiaoIZxmLOTcnWAxVeK
1Elb+lNkHRVIr8xrZe9c5Las/5HnRPFjdQ2xrNU/ggfYldAYKWLCgfD0ojCIDM3p
b8Y5/KFfqSH3ZcZeWcracuMtWcvXnjKc+9ByOFXIgu+OR8Z0gHrmp1ImXAWOF2PN
HGh/c/xlPtE1LIOscZFWYZbFOMG4Vs/zG0MTwM8Fr6c3AmP6ihbdTOKGxZTWyRC7
7OwpdOftMMo+1X2g+CiAKgrgtTRuTh8sTB9udmv2HXedt8W2lAKnrhDdn+t13+aE
5NZF3+c5HTau+GMnu6+71Z+NL+7IoTCLZ/Sns31NYtd5X5HxWkPPWLJFkjOrp9lT
dQCm4VV2Afe9r6gG7FEQS7LJM1jQ///61xoeaBRyaWTUrnygTOKicypURyxkJqmY
yHL+J681ZvHHkR31DxWwT4jK1i4Z9Xh9X4ue3p9jx7PXPzRwpQYbu1wxOAqUgokP
5wCsjX/qrCTXEaUhONVRJNj6d/iHNmwBzpavjg2x9fIDcfvOrBJF4B5YzlZ8wrQz
vwT23EdY4N7xo/Sz5e/w0O9aU+eeZjyh9/sc8zRsZXufArar/doWTaKKH/wjPXee
Cy4evzQGz8ufaX6eR8wQcacPBL4r9zbSXC/9jazZyUjc3OQsGg9po8RUbW6KJxQX
Ah384Ga6BKVwOJu9klVsRqzRLd1aAw8FpYfUm71LEhYDUJEzqW4R1Xtpv2ctb6Yx
TXed8SRBYOpdqOx30Yu+U/mkaNTmHE0CmHDEv7oElv/y/v978OyuT7OPSCncImMq
kVbAlGT9KUcE1/RmyJ8OYeleljfX8Pom2jOgBZsznvkDZOMJ1GO3+ap+K8HS0ETy
O16A8aMQlI3FdpiaXokarNqEMJfOJUjvgPAHht68zjvV65a5a1RtA3IiOlffafx9
0sI0GTK75mEijh1lYRHvzsoVYRzjKJ14rndq7+GdwRDz3o0K+C9MwgniEU2qKk+w
3dI8FGnKPBlqMGvL/7Wd4AHQVtEtH+/HMmNmoKtEu/hjyjZ07axzIWF5iCaXPuv3
TbPlw3/PICV+9aKWfrL0U2GppCsd2vWXwr0ttOVITqZQDUXh2QC1gmydMVtg6MTZ
e6ROtj34Rtr7ddltretf/MjPTPNrlUOU06QOpUHrs9AM2kcI5GOz2OiHmtTZ5rsz
8spJeOB+y3RlnVz7k4tFECU7ccsWFdW3gC/pBCopvY/1+2Swf1uJXAfMlktNOBul
dkCIh7kXCTDYgXCkgxHeCXpY9Zr+a0E4pa28B+m5Hq1tb7Ey7uVlZ/PNeJkd7VmD
ztVXLyN0YZGQfx8qKfDRcVHlbNGnirHatNwdMamhjqnIdQwC3ToGDdHFQM898xN8
Cl+oCORKIN2sce2aarlHtlaZKWz7TdTU4DssQNYO4pINstjb7ERg9ceOGSmThxCL
xcYiSKy/nPviB7Pcm9UdqDGOCkY3XGduocyyrEOEDFYeKd9grh4NocivpNS+QMq+
72AtKwCKdJID9eokD1OxNAxNOZeONJGa0ih9kyirDKhC4eXkiUbF5rum9319Z3lV
SupA27Wm+LM0pMWffQaOfAhFSDxHS/iHNEScr2w5exVFW7ZMkBVKEuU9BvQsuH6t
VFvuxsWLG6SQob+/14fLBm22AbE15FQvgrjN4/jBFDxTkKmHCfMmx8/lLNw4kPdG
pdtWnbdf4iosvKe20pjvPT9uFzxVqfNebGbzCaqMeALinL65nuy0X8lfkuUFeMuO
6Ol5gQjMt7QQzecg9tKtr47jebQ/Gqs6KN0ZDaUUCykbSDMNwg9uORpXsejhUuv2
NANfP97Gv2SUhJpa4XKIuIZrP3VlhM7iaolbN72Ky92fl+bWiT7uhjlKBhYfzDKc
VL4zaeSg0tYHE30zw+Lq9lLVk17xf+r/MJX8H2KgpQaGbwrOe5MOD80yjcQlk1/7
a2CDSgyZdbK6LgQNKumvmDFQ78E2/HxCHQUnFWqRyAsKSRsZaSCti+VQ5xe27Udp
plInYSHLp/f8YPCU2R/WzrhmTB8XTUm63n9bUOButkoczySh5GLc8ufN3Q7JPp9D
seV9OqSk8oyjH9eeTI4Nh+OwtTq/gsXgGtSCuAKMt5x5rod5LxAwmtgf3LESPln4
LKFeNFAZ+11uO3NZJ9m+taAbUMsljIHTccSpBQinvtR0c5lCJmqV23TsQQBufMN3
z2YDUjWmjXCvDcDmy4ee46mD+LOZTctDFwYjNEJC8TW37muYby6vPLdfhsn4xuVs
AttRx9sqbUKys3tUZOZKkkLKrZCMabUp1lPrMGtZH41o8XTug5hwmYSJju12+hsz
dcGheWHCjR9AeoUX38BjrW1OwQ9EZYyhiMyss0l+F6sxT2oz1KRD55a1d951wGWT
eCbzmaJ+RxL82/9C1FVw0OT88H3ChZh+jYA34N+w8sjYKJQGcfkkHsTwT6N65NNR
KuK74Q4ITSLDEinGa2UdneyHHomDIYMmstp1efD4bYb29aK7GAyROLsl3D6UZNtp
d8q1lbMgrZ1TJnY8Zl1MGwBkfc1XN8i8zyj0+NhUZKqQhXRsEGDrJ01yz2R2KCrO
GxGrLV6d0vdcr3zz+eRTaeZpAKKH1tlYU5oDeEaaFNfc2exkoIgK2ruYLg7+KtvL
3KvPuVAdtyS/yxMwFvxbEtjMRIRzBRelH2k0dJ1fEX4qZPKcrvkAvkO8cxIV6Tm3
DdwAiKiZXKi52eud/3B22RAGc5hKOdyZBbhDAeWYGlA4ShPa00RVIWkIs1oLELli
4yvFGPpZaZCOdrRVemxJ3t1O8X+UuGBICrKQW9qFHurUTR8jKlXmeRLV6eo1rtqd
U6kdobZLig3drMz1XSnBlkXSm2keIZ6uNXNmMMF//8RzJWwuMVJgpmqMoSL3mc79
dAA1q4bWJaaU+gmUiZbWS52Tpuhjh5fTx4tvt6k9ksz2PJdIx25kotHICAvzq6cl
Jpjf0bxqeZWa0kswr1NzbKzFJYaSxgJXELNuQNetWVp7B10fVZWlWjIH5oqh2m4w
TmvLIVqXmb0525AHVOLzheUDiOMUtw7ajl7N7Dg0manV0V+7mLEwcRzULx44eXYZ
4IC0de6DTIwfpSH9EOsMZx73bBOsAY0PTBja5dgMdUtUZBmSwSXM1qJVlSlW6NeN
dP5k5U6BR+wmCklgS+/rffsRvnDg1mbGCNFSXjyJzDi2PzIlLXKQNcAqMQ7dl0Uh
I4fluc2snaFHqq+z3Swefcw8v71i4kH465O/CmridlfiUr7iDXVW055zru4Usitz
FA44OHlcWIj6g6RQcs/ChmZx/2DWXMz32HtHuhO/gvs63FFINDqzzJnU3yKlLa53
vZ9Km6lfmc+UL1KrB223R80+ymBscyI+pW3LEZgNt10HER+0d6JpXL+Qej59a4us
2FCfrJQ/z4AJOoYWouXZ+VJIovvd0p0Ld+Fo07H8DgjZlY9pN3JDmOvBmEZYBayX
U6SKcFyTqlpiE/B56hy8gzwVFnewuxB9/F9F29i/xqltZC3Evnp4wk/6t6qc8Nlm
28N8uWrCtc01W7RxNhunbwxvCHYWu2zQ288jLLNuOYzpv5havabJ7go3+HBzlCm2
duiGr95TILdXDyV5mnt+m4c5T9Bq/w4z7hxXLk2q1WFGkx7RtETwGuqx4ijC8FAF
O5DzZRigAhd1/g21+ZsuSSmhGKBSn2sg7FGBL8M5sSPp5+lcIQm25a75dYygbRL7
mD/kyhMi/nADs5TsU1stdSJ6XzqGD4etxCF4siNSgH0VjXf0H0z8hQN8jwGnI/8u
Tou7WoeHFhjF/t+BvhaVQ0Kh+zI7EQPwgY+OgAgZSy08Nst2WadFlZ5+pYbN1PyM
ZjA93EGms5b/TYlz8EUNMdc4HPGvQumqci5Ii2630TGVd+pmmIIg6PGh7bXnt299
8rmBA4tHPsIn35sXUjU3gB+mxVFnpXRmEMs7r358w510NZe3DSuSISSl6SrsfBRT
aU1TfW6FKwNd1wE2F90uFYatft3zjRMq4YFcrV4m63ZBPgoxhkc2j+sq0Q+RdYqU
3n204tPl/JszibdHHattDiSKP3xeArjZ0WlnIH1+lRejaZ98fW3h9iKSfk9ADswS
t9cEt4e++zKgJQ2gZZyRAzJDC9QD8BMduXsCKT+sI//noYP9WFPRWjHiuez/gkYH
Hu9NR9PhIVeH3GZt6ZprxYtpbZUI6ZuzvCdFNcNuYU4kTCA5onHn10l2aOeUa4Cf
r4a2M3Gka7u7hNCdsM/cedZAEtG/LBD0tUrf6R4LxdcwlwFenjwMO3sUFD9nSZ9G
2l1ULyl+xQuQoC9VreVIsKcZfNohAsj8KvxKMKM3pO22hz73JinJLYvEZV6vRznv
LkkoPw+TVOHjeac6GwswtDmJufONyr27X8gJLHuDsLHgWClLjunPBlLmD984dsu9
8iZHqfD8WIirO2jYeCtYGOBKP8ZkeYa0mlScqfZ7/xlB3J6KOr1Xaf606T6caF/q
EumA5JyIuA70jHFy+ghNqL0pU5l5y2FlfkDkFxJSPQjl18S1/ySLSKNriDhFR2Jr
NWe+73MWDoMojT1N5Nt5HV6nLj1muh+arEBEQL5qbjU/qkOkYXQnYJSZXT5faHT5
Hcl0/etvJe6xwphWk/zWXylEUSoUidctR3K3DOKfevbvC915oJPi6c6WZNsKxEXm
bKzIGOEEXXCuNqrOzF/dS/Gy1ur3aE91J96Ae+HJkr8qMv0Amh1NR8fGrZsy9Zhg
f4QdcF40SYxth7JYKEnxg8hyALBXC9ubS2rv0jVHJeO6EoaDQI1rpA+W1tP2hxyO
HFTWfasYeVqG6CTm4ZdN692ry24gXxFEpmfRzY/UNUuQZmc9lZ1RYAXT8mqvlv1u
GQqKB8rc9D4Ut1jnHGWQaVmKfMl9CFYcQfpWHyf7hok=
`pragma protect end_protected
