// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H7S&0D558ZBC5X4(A,6CUA& )@/5M7N\/!>3P^*>9U!_#T0-Z.AW$=0  
HCB]:,P#UE V'5R>+5MM].\5$+^BN!]?!:M$MX\G]@P[<1-W%0RA+<P  
H>T*A8^9F73I1COUR5,$F<#;80,R92.=7_J^J.GA!XGU9F7VE4IL<(@  
H"R"88Y8K-90W*3W8"Y?[]@%P9R24 3B^$ NU!K6X=MIQK !$0>=ZW@  
HMJL;4R]RTH@V6ODQVI/5\T!VY:4#Y!N[OKIHV-D(8B'3TE(M)\4MVP  
`pragma protect encoding=(enctype="uuencode",bytes=6464        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@5:6^07<KBDAN(</2,7DAU='.@.Y*4L-7Q%^6MGD#PN( 
@JW\S,7NK@C5.TM2L*8BG_\$"FO$XJ6 C"Y[$&^;C0E$ 
@ALU#>@MH571V%UO;7OK=]CDS4$(1::/R1(# YVI.AO@ 
@M*4G07$!2<(WZ*S]W?V:Y9B\F9^[PHMRY>0;&0VJCC0 
@:JZ]!#,5-IT%5PG!<!FJQ2$US>"O5OH('.&JL_+2$(L 
@V3[YP+0?C/>7[%QA5B<CT Z6>LW6E;Q^BLEA16"GDVX 
@WNS26_F$WS+X3+"1&0FM;I@'1'_FUAQJZ)$RKCF2*PH 
@(,:UB#?0MIJ>OTN,-P_R*BQ_D8T4N+4WQ.WQ*4J^NS< 
@W= "<^%,7>DQV\!"[58JPNAM?XAY@9N0?<0(WCI!0*8 
@/1N4 3U1JZ9S;CX*MS6VTW<("Q+]^?TZ/N;K<B"04V4 
@6E*O]87\Q\B\\5U4=_&LOD,+CT!=71W3(L]J.MK^>\H 
@5M8J_>92POY@VOF+G&XR0DV%;U]L7"P.U^0-&;#6!<L 
@XZ&,NA-[*%98R8]3."&#Q=1X#^E"7>WQ 4(G2CR@LQX 
@58FW?Q2QO.<PY>"R*#=B %I(;1]NIQ\Y;%',7UV\ 0X 
@GUH\)*L*3<G-UD-& =+?WOU@#]/&8ZS4$ W'W'< \08 
@G]&$C*2J62-WP\"X %8/.')E27)E6)A5$,7D11<;.<H 
@EH7,H#7[YL7(N]!Z5O5K>SNF.SX4&:2]DU266HT'@<@ 
@#,;[AW-#+&;NI)L()%)\:%4S2^/@CU*25ZI0YG5SHD  
@<?G+XF'A8S-9.ZB*.QK"R\9B85=YB#HP,.\;"D&T0F, 
@*_[+\J-)_F8V@,I9R*WWYBEN:&NA79V"I"ODNSY=@$4 
@R%H2_P SO;_MG*4TJDX%F0%[#EN3D$J3$5^>JT:\%?T 
@ZJ#MF<"V>=R[W@W8E5ZO)]BD$ZN'$]9J*-8\#BT\Q<$ 
@';BH//X#B!S<V^$"\SY\9/-#-0&Y(_W/$I!$ ..=-:P 
@&_\',I+_U+W<,($IA6.63[L%Z?NM?9><'OOK"_M'$-4 
@&;$%)XQ39M$,6*VD(K\B\N)E" 'O1K8 N^NB+("5B3$ 
@JZ_:#+!3#G,(<!R6[H0>%2DCH==4#PUR[>+0X*#V0/, 
@:7'E^/3A96#R!$^DN6W@A/Q$C,)Z-[1\'IE_(K_QR T 
@DR2%5Q"(#_E ^-FG-!>F:<0)/Y-?+JQ<)3_T(;@*!8T 
@C@ANDMDRF:$EG[\G?PM<CV!6!!\]W G$/XSP:QCCZ+( 
@/4U4F/M:)*>6HL='MB%#^U!EE,:,)R45;#A;TK"G#LX 
@ZY!>I(SDO*/F4F>M/G_^F1AO$^G5] [!!"_22R69H68 
@R*]ITHXI5(A0%*T,W>?6GOF!=F A*\&Z<K)%D[Z\BV, 
@/L&M\A>:C-\G?XXT$_M"1G&40KVW>W\!:=XXDSG^MXX 
@Y:BN&Z'VA68"6$?:S4>FP=_WKP+V3'/]A.\F(R7A;^D 
@$CDCAA\ ^H!UFNX+::&A""%,QI#%*MY,CR*"7S@4"Y0 
@B==9)+&;YUN@'*L?5!2\75T:LEED2AUC0FELFD-8RY< 
@-(D"/C4$,;E[,8NBPKIU"Z%+VYD)J+5N&@@"/WI\D5D 
@@+6XX_T+PZNKB6S!J%0U3VD[AL"ZM89$^O8),2G_:1@ 
@-OR#42G-\Y(9_>9H'EF/G5([>T0D-1;K788_(*!(+B$ 
@PFLC<K!(\<V_U9#[=A4$J"!NHS*$N&6$HU;^-9QJ-V0 
@A8^"Q*TJ!H)O.7V29;Z<VVBU85]KU78YIC)$E<&,"Q8 
@6Z.=KHFEZ>SA^7B7(WT:2.!FEA\Y\AC<IQF\JO/1AY, 
@?2C^$VB/6O]9?.CHU<XCN_$2\;A[UW0X_()[1(0KF>X 
@H*G*F\Y;+X$,?(IR+;%T,16]3H^/Q(;-=\)!:[B51U  
@ WS]Q5_**[7TQ0R/M#Q2>:>)& 6AIS1T[-?LM[2K40\ 
@M"2;TXD+7BL&G5]_B>FC?K9V_-G>$]3ZNB]/IU1#61< 
@7_1%UE%27TRJT>O;WCM=T+^%BW?OXF+R+11'/H%?O>4 
@\+X",IGD<6:RAHZ/21 :,0)Z6R 9!L$$BU9D.WF2X+H 
@G)JLLB0D(4P??B69 &&V SX/FJ<NL?1I)%IW#;KN0%$ 
@Z.GY*DBPU%\?74ZZ-V1=6^13-*<R!Y$TBK[+I@K0V?, 
@WX!7A,0C:\*RS!]C)I:?KM*7B6W&\I0P^X]DH.<W $X 
@3 NUZ##Y ?AS/8LYNJ"MD1HD1W5+69!;CW4[SF-6U&T 
@^G]1=G%']'JUC9(>;Y9&G:1/M]@>-;Q^:,2#DG@!V*L 
@6.X\FA8D"/\O=<J&"9]TVGBBU,7/&/+5V(&I7?L([UH 
@J?A(Q_Q->)[9*G  -!X)7&A>3[8=2^X?:&'$72&6QML 
@ '+U@M4QWZM5XC-^9X6R[&_%52LP$DT7:6PA;%FZF&( 
@2SBE_U3=P>4%<2DY!KD>P K^/4A.G0]98C(PE<6?M/H 
@?TV55-Z0#Q+6AK"PDD_!.C_\4"M[]#%2XO$)DZ[".)4 
@UVBH*ST-OSZK)M!),RX/AWC$-L%8NH [S&K9GES(T(H 
@8VIYMITV#Y3^2ZH'D?<.#XVS&[9^OE(S0N=O[U+L"O$ 
@7W O42!,0]OKQF=&:HFF)$__+%?LF.C8Q(?I<B6FO[\ 
@CI>5D#\^E\J#2=FQBNK0Q16'N)0LU,&1>UM4#DD=1/$ 
@#P=MR'>+)W]@'/? _F_?R1>4ZQ1\&.J"Q3C"?[&H=1  
@T:[@L$ZJK7(SI3[@(5TE*9'OS[1RT4\^>SHOF,]JL]@ 
@S037'?L NQZ1@0<O9%JXZY#4_S"RV_R4SDH)MB*P&*( 
@!LKNF5W4<]2DGCL:J?C4'1/PPT%334CJ-MKK%31@>"T 
@HJ&6:N0H.8K*)@AY=@.\3PXAZUY^K-O &[ZL;K\W)QP 
@&[;G.)GNBZ*=.M^)'P_ED/F;M%V^$=J7YT[$-XT+A*  
@:JU]M1BI<F# S &<:54)?($S@;/R)?32-MYU*^C+V2\ 
@EQ(@UU=JK;ED#3Y97Z>V06_3>1K4###HJ$P]BWS[N.8 
@11&_:Y-FZ4*_SN3QABH\IG!^7M8[HV78TW7EXDE.MWD 
@#W[<74'P$DK'K4^=;8KXOH!HH AU>+K,V"^V5S;LGXT 
@=2^-#FM;I=>.CTM.YMU+*ME'-/Z0?ZAU[4PT7WPEQO$ 
@)N,G&V<11M-)PH_\>96:R""A$"U#EA,?UPE"G3>?%4\ 
@K<IRAG-HQ)*]/&XL@)7]^(TP-]$&2" *-L%HJI3,/.\ 
@K=ME5-J?)$8&O>RRWU&M6+G]2>]E+^F=.1'V"86P5SP 
@OH3,2',4- &>?ULH;VP="_<M14$T2G8$TJE%\).@) D 
@3;NI=9B N_]HW_=RT%RXC9ASA-7.HPT&'Q"1PGF@9NT 
@":!@CJNY3K^8Q_8.7L.VE53?MR"04FC-ZPN\$CK ..0 
@4@2(3"B;XQ=UAPR!(M;5D!Z\U@\0]ZK+ZJ2R+)'T59, 
@RPM69J=C!1GQ:+,;F'K$V0$8WA>D=8CDZP&#7U\%Q_D 
@B,*+<V!!.&4A'H:\>0LJ;=Z0+C;VI'%;VJ9G$K"XYZH 
@#/@H%K%2"7JM2$C6MP]KE_3O+6*8&OS^JP(VI,<H._D 
@Q*6I*ZW1><GOVBVYB9\IS1"NE,;EWB"OXFF2BWG[=+( 
@S.H.$[)84C3KM\25194?:="HTC&U,L*YDD$H>AYNH(, 
@2G$UH!1VS5JTDPPZ]JUF-6VOR#X8 <3NR1%<)AP%#Z< 
@M#?K86$Q!DGO%,Q%NBJ%.%_P*[)$<4"S7+6&C3-?1PL 
@'@@37).9KB8#\:07&EL+++IW=#B(=48>P*HN+5Z^'5$ 
@*"FIEF8A/1:\W%QG=)\U(!U[ ]0U&*.UF[-O"K<S%&X 
@5S;_,S? O!7PT345O-X7(&O((*H,75 [[IPRQQ#MK 0 
@<&TN#!X?]+=^!8^8R0U3%'9=;5Q$VT,NYW_2NM7/O%@ 
@RCN%9@KGZ-^.X9TZ)W<_PI[9#@]R&_&C;9 B8O%6Y=  
@\A&\" 5?6>R7RD$E_Y";(_MR%[:A(B*.QG^8B"-.P'\ 
@H'>?*Q(AMYRA7;3S:H5MCN05_=T1\[C[V4#7&[=K9/D 
@10I=J4T2J@.?88WNFH/VAE;,]9W'5,F\N,82!0XV-?, 
@ZT.?;#0,^L1TL>J?TH1.C'T1OJ0EJY)2GAM]@QKZG*L 
@CG7AF@_BH+5+8N3'2.<Y'J_-EO/9VG2($-5/]E;VJ%D 
@6L;)),=(9XQP^]@,&XK4EY<5#4X@G&N)Z(.54YYP1,\ 
@!'_B6.=,Y)E(U6F$_X?H% #Q[#T0XXO_%CJ4D,XYXJ4 
@UQ:\"K)%^=I>>V;6_J'CKY.JRZ"(3ZI[B0C!@5 )NQX 
@G]_EPTS$59&DJTWS%+I<QAISW:J-8VLZ/7I!DKI13"\ 
@'X#O]&ZN7<&CH8!9_#^9$BF6)IJI;52CBIKZR:8Q1KX 
@KK>!A<*8]1I]<J2- 3;Q/GKF"4^:X<L1RKE!V$842;( 
@-+R[F:8P78YK,OZ \BEO7Y[MT9:4#F6G?'?@Q*C6E*4 
@]X[Q5?J N;S!)5<(%:)P')8Q*,@L%$;-A\]<4'O9;24 
@V:/Z:WX*_-Q VCE*4W"DL@]_N\JPKS'@_6?C1XB^D9X 
@7P+]1!$B\E.XSH&VP4G42( %J2]'P;YRR-A^YZ]9-EH 
@B6U/:_?Q\*\ /0FT&_)U)E#3^%-_B)*8["9T>[;#M_H 
@08.'%-U'3)Q7Q^?T9*I&U17X3J8#>X[E7(IJ+WDY_,@ 
@7 =J7FD219S\"EI[)GSP<U#;3;1EP.7KUWCP?0R-XHP 
@&!-S('H;0>\Y-!53YFX.AYIOI[:63WHZ<P/1<W9#$"@ 
@OA%G(_,WKCZC.>>[&0&*[ J]\KV/I(7'3<;TK8^W^UH 
@&$(OYW9JQX,0J4PK5[WI'3@O0]]JI85DK6H9;@'MB8P 
@V3@][D1-YF@NT8$FC"ZLER0C! .^E@+\)I5C8?S'G]8 
@[$+OW'$,])5&.3'3=BN;C ,:P%]6BLW,ZJ^LR)B[;%0 
@Q&DDMJW8BFU!4T+J\$)PLSF\_VZ8.7ZA:Q*#_F<;I8L 
@FTBZ2]C6]@1D@?J@KN_?"]P<T9G1U"O^](0;>M*\W>< 
@XU<VAY!)LB28&W6YPY>JL*S?DP0/$V!_ASW?.M>P6P0 
@T]E #$YLHG939J8DXN![?<+WAY)249KWPN9,^6DF;!, 
@US1P5+XA3#K*5K@R'_)2@16K_DJ3,O_8 ;XJ;@4XF?T 
@,?'N.WOH(V5/\.K.TL#+@'VM? M>%D;@KTK!*].3=]\ 
@K1,I_/$N;4D8R"[+\0=-^@!.3NAL/%5FFW1,7M5Q%7( 
@Y<.D4#P7E=.1M:_%-A%&%UB\3Y^)?*4 \$HT(E57!"P 
@G[M(KFJ.=,1V:@M5E4V4;9P W,E%/Y(N]@K-LDL[CCP 
@R*,!89]EY "!CV4[SWJV^62U40;RK2;J*#Y;F'B<-M  
@Z9:63[N&[74\X[ +X)*L0";PW )0-*0Z=BK8JL*A%3L 
@I0$;HU IT?XYJ@\1.+\D<I;L->TC.Q2?4! M+F[B'V< 
@05YR,\=F[,AV*3S^N;Q*(4\(E74WA)DGU;I)3JWZ5,T 
@90U7_ BT$.2NJ!/4'PS/D9K%1@^2U@O*S20<I#</-2H 
@ZSA<"T("NGAQ,=CPSISNN?@]T,YONZ!91U,TOY$WG28 
@VU\9- 7H;3GVP$W2')N(XM5Q7PBF#]53=:_!A6XS;L4 
@E3)Z[*2!%*8%HN/'Q-!UM;-Q3[95&OF$RK:]026.2&  
@-3 U3=A([=E(+@H=+WZ)A"\,?)-4?\1'[Z"2I38V")H 
@.3/"W!9P3!T(;*&PM1Q(B(DY$\ UH2GMR&&)UUV/Q#0 
@YCK8_T@<N00H@=FP Q!$K47BTY@D]#]DV_G,B<;#*^X 
@YQ]\/K>Y$=(-*(2]D5<KN*'K!\B^W*"IN#OO9=:\M34 
@);W]<AJ]?I4C^Z.D",TXDMK 8//\G1C#AQVUOYAK.VL 
@'ENX087)[.N_@!TV[EV:NJX&0J0GODL>8_B'7B0T7%H 
@FRRF=A_U)/RO-$9(5X@U5VV5OE=O(FF,PDQ^8C)-EJ0 
@,:T;YL9>$UE'RWQ;U:+"+4FMFP<K.69H*W?TM\0 (CT 
@?+C_BZKY TQ?WY)40?P5;"SZMX9QUI<2*\>T5HBU)O$ 
@LX(HNR #E;A#+L+HZ@LW&"$BEE/#]>\ZBJV"7X-8VB( 
@.L^Z<S(D[OT%/11$RT!)HRF=K\O1#^K RZEN1ARX=#8 
@?#=]65[[JN19 @9MENN6O->X#_ NKM5QI?S(66N>4=T 
@JD1ET3/%@I$]G\%?!2PQ'MG=_2OD#PGDSQ[6I@WIXG@ 
@&>.!UY)5KZL/?EM_%\E6<9^ 4)FK-S[3;SSNA+L[1V@ 
@FN_6C]4% R<_77LC_[>+M<#N)7)9W%30:<)Q4!9?/%0 
@$0NGW?.QMQA7@6*A?"HQ?Q#U@TN-CK%=&=97=[_VE.\ 
@J82.2MVK6[K;_K+Z2=:ZT(] >F5'?_/#:8A"J?TW/:, 
@H-C@KW(V)_9;(HN\0A'<5M*<"] ??[NG,'#VU:GO;R@ 
@N]2COQDP#O(N#O$6_NOL?<5CHH<UO3V[3UP>_&'68(( 
@P%[X6#.ZE;H$,Q9?4XK&I3O0DO@H63AN[+PH0 CT&=D 
@/\7N0$<!!FL3VU+)P>E=\?GP;S><@K'(W)3/Y<R(Z&\ 
@-LFE_Z<26!J;=\X#PIX4@IJS<.!(AYHH%F&CS THU[L 
@%L 13/O!V0("]2-, HTTZCQJ6T@DN(_6P%B#$(VU2\0 
@#H+2.I1-W#-2Q$45LMT/_1N1EP*BOFGR,+H-4_V .V, 
@A%.P$A?H\4L"08SO<A_-&S69(WRCV0K0#JFLD_X+6B  
@E'.9Z&+O<GZ'9?;#UZD.=L@X+9TSOXF@@L^Y+F[FT-H 
@Z+K-8#7MW&6S3PDLJ=-4O?\ON\_:HSFB=5Q[9K+"A[P 
@>KL6Y'WZ[&>#0TY>^[PV_2(J-V@IH%Z[::V7MC1/[ < 
@?L[.7$\E&V9ZNJ1:C,V*=^Y<E9N4;]>!C<(7'L=9 58 
@RLT3RSI)G.;HG:W%#PI\$G9QA#J8]3FLTN*C<QL0Y;, 
@LCT5=RLDTM&)B'Y,Y"&P$'=_%A+/F"^R#CT_(P'->T  
@<M=?*+M3NN]F[3L!$ 7$K$21NUB#8XT9\)L(58'JVQ8 
@.XETT5R<>*"N-A^H[_7VG(!]FJ/?DPI&QCPN??3*ZX, 
@)V-\-L^]8WB.TQJ ][*O7Q[IGW)6/(B$+BY&=3#WF:@ 
@ZD ,<T _D_2;[4!9)Y9A8,6FJ+>I?+>Y*#&+ABPG^Z@ 
@3,!/QXT'^A7-H)J^L0)E=?&FV@K?X1<5!!)9_[K\?-< 
@JEFNT_0BV(Q*OZ*9+E].8K)!1\#19Z%DVC@.?V%O7R8 
@4A/5P6P&"*J%'>XP:3K2#L:&YI%X83S]0%>[B.._1$, 
@CJ[00P_]@)Y!Z.%Z"@:7& C-NCQZ&25YJVPC<E4ATOT 
@V57?/EUJI5-G9 _EU6L*HV]QLH?@"'P] KF))Q%B1B, 
@/3JUN:#W4N,Q5/M;.U:0O*K"=X1O"1A7?!MSE5ZDX'\ 
@A(L;E=2XYSU6GVIK 5&#A3:^\,1S+I)'5U_LAOB]A0T 
@I27EXR^/*JR9'LS$4\3;HVYI04&!21E\VGZJK!*[;:, 
@K>O+/9QCLBA&"JN,00]Q;81MLLZ=JW4,K&E7<ST9\0  
@-O*;KQ9\[%PU8*_L29D#J@"<FXG+]H<FF7TE;!YES3< 
@XV97_Z5G7;P ?W.M11)6F7JNM/'!F+=Y_3V51T\!O'$ 
@L (@Y]#+R[#6V KM%21Q>OV_O>QI;CAZR\TO;OF+%B4 
@)BI_WK'1@9) M;A >HU'RL::0LB/]:@.=L08)/I%#0< 
@,>@ =H?QB=7/,5S G_S+OV3>%_'1!1MD;X3SRA_JR]T 
@N'RG\W8))%&.S?T,Q0E*6N6OD&5'-W=RY2=HB2;BQ5H 
@<@RM)O=>YJ98P.B3(XR#R]H1/%XV"B&OW L(?("1^)( 
@D)B_)Y)164NV9WE"Y/?37DR]UA]7K5@?+#5)G?(BU:4 
@.YGTJWLQY%*,=FUYR3XSG=KBW_C77\-B,!2"&+ML7", 
@DRUQP]X3Y*//OB#8\#+P*8M29IFX.$+M;T2=B0B*LS< 
@_ .X/PB6=%LMG1^O8K9HM>#/MT$-WM:Y.FS);&.:UZ0 
@H- GS0<W&7M^_-M.?+Q['U0!F=5$/Q_;TP%6[Y$^S(( 
@E[WNI?VMR'8AL:LV8TSS[;E+FA&]"8$+_=M-^D4I&]L 
@G!!35<NZ,]8(+QP A1((.^G9']5Z0@C9U_["<?"_F'  
@>,M;#.H,A%@'(H'=*E(L5\LF[$'?Q&D*:/^(N-_$OP0 
@,:G  \VIU2J)T17(B"1(!%100,)HS)_2GN+0I)8E[+< 
@TF3$#L)%L).4S,J@VPB+FP83WUID03>8''X1:=AQBQL 
@7SU!K3D7\H/6?@L%R7]!2Y]HDHJ$#D>@M #=-^9T2/\ 
@4$%MI:K75Q6"T\]RNA).$R"/OY#5]^>*!QTZL*4!7=  
@45XT1]-WV50!+@'IS0[!TR$'?%M3<>0L9WO1B&[F)0< 
@%.^IU(TTV[_147P%$+E4Q<:D%BWL8%(&KVA=+ 5=P.  
@<ALZ?%XP<J8A.AQ5S,< F:A;T]1WKJ9W@B<6"5*K<^@ 
@UP'0KD]5#\->TWVFX3##]]\>5--_:2N\SYXP?NI^)V\ 
@_#^8#\_\KT(<2KO[&C E3LL =;X"KJ@S_;MXJ&HU$!, 
@ZNW$:@Y\WU-1SBKMFBYGO@!98/NLR6!T\TR;8@V*7V@ 
0_ALQ[K,X2T2><Z:_C' =[0  
0RZUJMNC8 CR((V@_ U/WK   
`pragma protect end_protected
