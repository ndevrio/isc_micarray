// cic_ii_0_example_design.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module cic_ii_0_example_design (
		input  wire [1:0]  core_av_st_in_error,          //  core_av_st_in.error
		input  wire        core_av_st_in_valid,          //               .valid
		output wire        core_av_st_in_ready,          //               .ready
		input  wire [8:0]  core_av_st_in_data,           //               .data
		output wire [18:0] core_av_st_out_data,          // core_av_st_out.data
		output wire [1:0]  core_av_st_out_error,         //               .error
		output wire        core_av_st_out_valid,         //               .valid
		input  wire        core_av_st_out_ready,         //               .ready
		output wire        core_av_st_out_startofpacket, //               .startofpacket
		output wire        core_av_st_out_endofpacket,   //               .endofpacket
		output wire [3:0]  core_av_st_out_channel,       //               .channel
		input  wire        core_clock_clk,               //     core_clock.clk
		input  wire        core_reset_reset_n            //     core_reset.reset_n
	);

	wire  [18:0] core_out_data; // port fragment

	cic_ii_0_example_design_core core (
		.clk               (core_clock_clk),               //     clock.clk
		.reset_n           (core_reset_reset_n),           //     reset.reset_n
		.in_error          (core_av_st_in_error),          //  av_st_in.error
		.in_valid          (core_av_st_in_valid),          //          .valid
		.in_ready          (core_av_st_in_ready),          //          .ready
		.in0_data          (core_av_st_in_data[8]),        //          .data
		.in1_data          (core_av_st_in_data[7]),        //          .data
		.in2_data          (core_av_st_in_data[6]),        //          .data
		.in3_data          (core_av_st_in_data[5]),        //          .data
		.in4_data          (core_av_st_in_data[4]),        //          .data
		.in5_data          (core_av_st_in_data[3]),        //          .data
		.in6_data          (core_av_st_in_data[2]),        //          .data
		.in7_data          (core_av_st_in_data[1]),        //          .data
		.in8_data          (core_av_st_in_data[0]),        //          .data
		.out_data          (core_out_data[18:0]),          // av_st_out.data
		.out_error         (core_av_st_out_error),         //          .error
		.out_valid         (core_av_st_out_valid),         //          .valid
		.out_ready         (core_av_st_out_ready),         //          .ready
		.out_startofpacket (core_av_st_out_startofpacket), //          .startofpacket
		.out_endofpacket   (core_av_st_out_endofpacket),   //          .endofpacket
		.out_channel       (core_av_st_out_channel),       //          .channel
		.clken             (1'b1)                          // (terminated)
	);

	assign core_av_st_out_data = { core_out_data[18:0] };

endmodule
