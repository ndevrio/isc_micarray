-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
BDWHU5cXD26soeLenBJNvpcD6bgtU/6d1tyOQ5FgmAOrzLxT0VY4pqKBNzmqkx5N
NI/0HmubczWUPOZ2IZx4Ad7f95b1BJYod/l9ET5sGKRn+nzI+maFqVziglbU200I
jcweHcbIWJJRfaAZvpUcnWKWLggiZ5X1OSmOA6aIdAObzNxAYM/a2w==
--pragma protect end_key_block
--pragma protect digest_block
sJelUufG80tepaFyXrbRGDF/GXA=
--pragma protect end_digest_block
--pragma protect data_block
Z6YRvXlTzDb6KmjNPD1zLN1w6/hLACVxKvFWLP2x+Er700YsWoUURwKcuYn45nvO
gEt1k3nsmiPaZxHzJHtYReah0URpojmPpwg/dLskkVRFuGGaQ45UVWCpMcOAQQTO
gY687yAYs7AnCzfGU1kc6p4klcVphgNVEs/AyowtffJWx1ut6hST1aAU04Ljk5pP
bCnAZeEo7bVWdiLotZfo82UBNrpMGBfye/PH3HNfxDYstxmxYDVYqAXAZPhlvrGq
Dp52eumArh8j75X6yjjdSps6c3yxofvLwjXS7QJ/4I2K7+1vriLs/FMk+yRN8Hsl
gIGLO79q9/LwG/oJdZmQqh1yMTjtfj8twD/S73SYz4pPFqIFRpPFYb13dETGKEue
X797putBa/XMG7TM7Ujw/6E102B/J9fFt8tnydiEj8332jx7Vrf3ourk/mGe+/hh
ro7vcNyWdMAksxvIBgI6m/L19Rl53RsoeVqCSy/AlqVw6p5YZJtfwjTCoLMXUSt3
2NMnmK77jvi/PWQf54rQy+1A1S+w7qvtWkWh6B4X6YqFCoL3Rh65g9NqXR8quOYK
rbolKdBItWy2eADEobzgKhqHCUvfY/hB83b4Is8oNBRLjHquhpeQFGdyGN7SenN5
0f3ft0NSvVxpr74mBfy22F3YkwQ1Zj4d4blvfNFso/gocZLrP3LJ723z6mQTIp9S
0tF4LVAkyWBPU8IKYnvy/YWV62oNrHmt8fgZIbyjAKEnC8bNcypzpLeSmw4Lr/y6
d4/2a42j7QjDhEqXvPwUr52B8hCXj3aERTpnZMVaffYefYIrax8aRkS7G0/RIxzx
mEXs02O0qkL8pAQ3H9wWF0N71vtKVJkwcykuysqD8qa335WPSWtAVjXY5xwreD3J
OVPuy73rthfqB5nkx9MUdH5HwWHYNfB6iSBEzf+pqetsLQF8U67uYb+dbQ6qwpYo
G6rNp9sT+WxkT2wTWHxU5oHoWXYc86p3sG6bu0R9o2K79ho7X0H3ng+6U3BMOB2z
egRMnXljzwxBuphnGElTdfuby14w/6/7pv0dOCiMW2R655761KA0ebUsnZltu4F/
rQpej2au/Ne90UqeKd+AlKJHgC7GCKDdypw2CgH3xORPVnP5irPhyNWdFG78KbXZ
Qw6dFLDFYve72VFqmh44Un5iB/UyBfnVe/Up0Gsg4ydREZiFTcMnNyw6pXJoPHGP
o2RlN5f9k+0kKVd4F6j/Jv2jxJyo5Gwfdd+g4LEf0N6+RIxwST/a4CKvVwItC6M4
ReIx6/6IgM+V/aoKkcWIldkkyXmeEx3Z/BYZWlLX3zLWAQ452gC3QyV+q1EZ5Ix3
Chmno61KwgqnwJltDRE8rQl9X6DaYQvtgS9GAxxmjWxoIwOOzny2du+Kc9r4vGhA
TgZMaVT1HQZZA0VNALrwrH58rvoM/AQALkmRkkNmNaBmvy3+wqBiT0uYxuHQEBjm
UYIjqM49VgZsHcHvfayPW3KH+Kt3n6GhnjJNxYYf32RxQ4heLlpTMtf5BI1xTxqZ
uTT4b1vU2X4/9cbIRFfgRBLd50gRD5pqwz81LMd8upLKUVHicWQXshaPTJOgKfC5
YfkFuxDdvdZ1D4wzSkTEaC5BamyIb8bO7VEd/ZaOqwp/I6MC0NG4j1UdnMyxlt8Z
TEzYx3hVatzA8UzF4roZ47UlfUpH9ZDW1FNzr9GiG4xT0JxSSuc1bdMFdy7/ivdz
W+W9eVB3xDTB8CF9RV3lgZZigZ0SlgH+QfeNR7epbSYr6fxrOyCMW9DYrR4A9REC
3PnqDSkWoe1GxV/FP3gWv4aca2HjJEZpiZwv53j995NCCtL8shDXjUdrVELg3EHB
rdDKKU+2t+lzS1Q4n1soctqKdgtBQdnr7I1XTRjCNor6fwUUI+cs3Q1h2DNdHTjd
Rvq/i01JShBx5MKIVsym4kHp7ZKixuO4xMpuDLakUeu8/ahVcbTUQnDkFS9OuFBu
tUpoxsOisksz9GR537bihRdB913NLCDkBwqAcuH35YhoFau6bqrFX5GK+YwaUo1B
TXFQ9W8BdsEprm1G/rAwpfs6P1AfOLdo9ecnxMmVoz03i3Oep59kM6aFSaWMT6OY
a6nUVXQvKBHiV2qdX8yMYYQi2FPHRK5d45/9EXV2Jb4OzoyZXsvVyfqyiPrghOlt
M5LTHmRgq3ChKy2LSQC1aC5qp+OiU+3DR2CIyYd8WxijarZ9UEXcprqCTWiFnRgC
h1BQEP5gFktKtkbr6Wyh4g/vQ0SnyWmOGZSSk0+Ttj9/xDSU4hjNbwHG8DvOKawn
X7dICEsHxnJuhbq9E/rFOc6K1RyBT3lWLF0XyJX27U0l9ZeOROI9IrPECnCfrEL6
CF2gBQgfAjMA7pd+BMmIXWKTaHCX5QeQSpBFzv8w5Hhy3FHxhPY8xw/7sJGFuCV5
Hkx+tojGLVvQ6ypsdIpFnC0o6HTZaI0CcOxQE80D/njTBmHiBHzET22vOsP+g8gh
fg0adAclYNOGgxfuwfRHNSjsFIinZHQq0Juy6w7sv4qnjgG8ADlto54wS1VuVQwD
8pvtynTgZ3rbDZVYJIpyENtt1hd9iFUk2h87xPq5ak/wAftLiu22BZJhA4cJ23qh
28ik8RInBsVifFta0gJXMSTXDL0U8Vk/o8DOibESp3p1OXXP/P29xiNkCcjEW+a9
2tCDUISgkHhtZyvo5YwyRKFLcd3UDf8Ho65rhoe/TFi0gIfxtdcwjxVlucrGZjzC
D64ifwS3i/HQ3KyqhcKfvQ9cNez8ApTxULifXLnmbh6tpSkjy6jrHIuQpnoI1ZUo
2ijQS91UYCZ2qRMkt33jj3oYnOFjiq0iJKk9F8fE4Zqid+6Xhshp+GdziUX3Ou05
Uoc99dLmskTs47zA7Xuy7uwe68KZWK9w8ZTL1nYYwd0YpArCE6J0xXdF8+4fx4u3
7sm7uWWY4dia+v4NzODyhPiiO+Mqym/1lrDlRpQ9IYqa1lfICrZpnz3MqANcFFE8
AzVHHNLVDAHg4XmdXk8LB6EPMwUpzmiKnG5qTD7IR0juorN/cm99iJeWYM5KzDCa
8pTZIODOZtafF4eON9CrgtqOepiYwAgN6gCNYAxbCEySYaOjuL0dR12oP1HxtQag
2eTQX70KUiwZC2oWf0LguLi5+YksTW5/K8TsFT+La/psSuib2bCS58bXuk6kgXlX
tz8hF3v/GKU8QxjzenIACgOMdFkYrTsJ+IenDNV4Kk+RHTXhSZbPcqOoIRKrHkth
ZT1dWhOfVyV2fzknw5Bt3gOSfNcKBObou9y9V4zViAx2zP1ASGb6eLUSySEQnt2u
znFxlQ+oNZYf/fdOjeqRqHx2VMLYSahv18Bv2uXcI0/zx9MYF2waVqgcUtPUdGO9
V28mx2PTOA7tP/YztO1sWnQtf44D+urFaQcKOuITtLuHoXh1Mp0W4xrpd5N34pqn
mkt8k6qWyZeVXc/CBUKz89BgJmJzETyMU96iFVrNl0xAgfJAMpwW77/TRuMazfxv
J0G+792vlFvYxWrQvIG4z5OzR8eGa79/wQLlP0cEygRnTX6gWuuLb+8ZBSPypPF9
fs2SwbkL3uq507fed+MgpgHJMBEs6BIPlD8w9VjHoQd36bPQholHz/qUGWC2cjzn
W9AXX984Un8RrKVveumWgAjpybZQTETkZBnna6okdyDS8xTJeYzYF5pyvczPGfFb
WjUtXpxaRWw+asVStH2XFWcqjQB+og9+fMoiQg7XMqQNd0dtUVzEAhZ0fyCyrwib
mPhXcH66btKoNZGoYeqWhKMO0+scjuj2+QIy88MlNsF6bsAFtIsu2S1KXPzVsSZJ
Iw0jsG+N22VYcP+4qYQzqLrjzNJMJuSHMiNd48oBIID9W0FextcL4PrpxSKodOXJ
iZAi7SOHymPEgfIqUrcb0k43Z7BXnx4yMz9/LtCCrAe9QPA4y19Y/pSa2qvTlpXp
YBNe7mkRnspCptmTgAo49gywxzYfcus7I8nOIvHvkjbtZLZ+yfMl/02BFTM/2PJW
sWrgu+7MxkjAU6uq/bOpapY+b9kAg8UgkeddpiDDJNeI7A65NFCJmv9WQUrRY0fy
gIPRynW2biyhvX0QR0qOkRx/bwweqB2M0OdLkUilsvJt8Pfi4Tn5jHTCuYUfslMn
8QO2UC101pE8nhgWrwBJSWFX9Mn7ywbn7tDVMvNPPBHdulGYpYrHPGVqzK5h+GjC
n/OJyInF5yilFL0GUgE7B365aheyW4euhhs8ltXJpzT2+2e45ZCxcdPwIDAWhf87
PRa1NC38xyjeTk+nacNXHUJH5mkyFRTK3CMyiT7DDSJREoUdCO62vIapJr3ri6pq
4Zf0UEa4rK3cRC7MVONC8DWUnarju8B0Ia4zrWxJSZXVGOHLY158/jonMqkaWjMn
p6SXjUsjlHZOawcj0z2JtAVbHOdfX30DkZkQQfZUt2uLPDeQNUFXjL3A+yrIcxMD
h/6vlw0ev2HmB1wh0DwkncsiZC96/F7UvtP2vW7NApDXbd/y+6QQVyYXZRYo95lI
Sn4KgEmbGXy0L7CXraRTWDVkn6WJBGzypUhmBtobOpQG5xAosd7tLbzKO5sErtDa
/ircbgKL4cnWmNUpNwr9Z3tQBoE33ZuTprL7+KheliN03zM2WRzWRgDyV4WUCVWU
FsafD5KpLfUBbKlZ6yOTrNR3FScPTPyFA9KGw42Q1cuePGI/FpsctFY9fHsIEHYT
gOOvl7pamSzEjFnMfTRqL0lcP4fd9y1ubZQXy9NL4Mx6K11sLoGw5a+tAYcnnAf4
tFUdVJRGPNBkA5nURArXFnq33qdTS59if7OMrZkhVVxyykyZITF1XezfY6APKXYP
bnACRdqByqq41DzHSXaULlj7LHJcClX65ZUhhmplawoDcPRko4jEuFDTFIwVAe1j
4HX2dAXDT86guXbn4KcbaZScT7Gl4ybb1SF69LKEQFBCqID/gqyaB6KczBvuPreo
Bu4gANjEncPYRNUw12CJwwRlG91NpGBp7xgm2lYkxRkyNlyALHbmM1/lJYFjqAca
ugIGZhjSWFeBaXiy4vsCvWcVnyzMeHkRjlKohcFEvTJfW3E4v2sMEnw+L0lS7tSH
VyHFZ9RRy1SLZiVnt2JiNMOa3AO2an0QIvR1X13rsrLun7N7PimNgbnotLM31HUB
xq645WebnzKdBHNbBoWpE5KhgbUCobuSR1QF875Ls6JNeIeJZ2FYOAX8nXGqgv7J
4Rq0BPdKiqV3V3ggTfWN0tt//RH1nL0mpmb2kRb/9p9f2W9cEQ0Uw1MzzVmMN9t6
Q+38y+CJXPZRKQt/Zm+EE9J/E6QZx3+zJOsAt4iSwXMLCP+6Evf1VMwrAeL07ytp
0xObAtTF5jr0eRjthx08MRPFEQCC0p3rKjlQrwBPdOxoK+4PlBUaGU5T3cFtSPVp
3XAMeSqf7Hnpxgql3dOzKo++uqMXUqCEDtdJ1Um9atgp/GVPXVcgeB+2uFkJW/pR
wwZZG47lgr2a74qERvR+DASX34uUTkXj9CmQL+wWGeD3DzBaJGFjr80wb1n71cX5
45BWVWrV65ymIHHxkFGHxmD5pfwaxIvCWCxdeR3owtwCkFLKU8zkFamzRP9iQlzP
71fjFdDllAXoWE0vDbvbVHIN7SR2Hg74Uk3XvqZHoCFq++kbX+36FNKm0Tbc9DVD
Ijw7mlBCx9ATr+Yw68n0PPkkh6XA0mlGFGF8i/rPTMfWpIHpJTRd6rXnMai86y8B
4U1HqSJ/IZdbrBJ54Iw7K3c8TjRSnHK5vRPMjIrRvlgMMo8GhpJoekyerNsT6uri
EsXnoI/TjKUEOje8Q/EPIaP33nn7G5sut8EsTenvaZHS4pTBrmUbm6UY/mrCZ+PV
1W4fZHx67wEqAlDT0egoIJN7frirhEpgblumoL8SPiyYgex/gIOd1Be10TNXgIUM
wVPOTIZBmHaayVLWnEG5fxo0EI5Wez3E5KHYy75enKIryx38drCvSBl5DMmswl4b
QTt3ssfrUOieo/VGUtTV29JR4kpjhlbSJzrYb0pVgWJ2QO8OjSgq9dT+Cqj2se7R
neLZMIcav62zvF3z/CyTWolccjN3swXMzO8YVE30XdLqy/NhCXm4OoPyOBmNzoV8
wtlhqiffDCU/3BzrP2gn4Tn5vNy+xaUZp6yCLW5mRm678WelvRXc0joReiKv7of3
i0qqVwV4qFj5UI2dnhkCfKRbHs+bKWbP64bcCZqJEaF6ly/9quvaB9qaKueIpbUn
W4p4ffNgFUI/y8ou6Gy3My9Jq7WYlY7gO6ISVIrLA0i8gUqJB4ctwdhaml9tUoS1
S0VvYDR8oKXjwPZ+xFj74sGckc1kAoTvtNRf9xiWrNbSu4tTKPH02l+XSyLFUV/w
GNr8gB9GsqKSkjd7AcgBRcgUNj++whG8VDLhKXpcbm3H1niNOmvvs4/acby3Btgp
4Mz3s8bs6HbnYn7r9HWvrw3d1lBaTYvFLvjgIlj6rVqUC0QHgZK9OXSmRwQzxW8n
oyWbnD5gvjBUZo24IpgJT5qTK9rQB/yLGJwOxkiYx+V0fEj3g6YBaSKScJuBdHB2
fFohaNoXr8yKkLSYBaHiEqLvqx9ehvEsKPnS2sEEA/kEra59QzR39w7nsSvlQlxZ
zFzlL1mR6/2WOFIXKR/OWXa5ZFGU0h4nYtit8ke4CLROjm34d07SbAxLWFW8szUJ
uyc1Qmvo0CfcQau/CIvyhKd6apbz1WW/ats0XezqK90s4lBFu6bVuVTGwyqCcSsG
BczHfEYnEhM+S6BeXFHLGQTRJN7FtCr+Ep9aAp5FZBDt2JONQ+usf+9schRZC04a
H4p2Ro9lZEqCvWXDHncSnUGbIN275QKat+Iia8TJFx+g2bB0BO5yfFlSPM5SCNUr
y1b3EnGlcnMbhKqSyGNeH4Y98WnUCQA6HhiExKv2Wm4rq3nidayoY2LShfy7RD0W
wspzxS1SMGwzAGdr437VyQu0ZdYG2++qog4+r7a72D6MAkFbuuDnnRLc65uPv5Nt
vvFTR+urVAFkM3soISc2vh9HEfu2thrcaM9IeN8NOL4qzTBPGcbX+h37ZOv7YsK6
eARs0U6TpnYLZzPJ1wjdVJkCDPZno5XizBcOEcPFf+i60/7X0ymdvUG/tpC8yeUN
FThosXejLpkpaiZNn6EFpV2eOD0blrw0KxQiN7yKUiRDax4omjsIlFrfjpzbTjPt

--pragma protect end_data_block
--pragma protect digest_block
oXxkz1C9oLQD8ZFRYNCJAVM2KyU=
--pragma protect end_digest_block
--pragma protect end_protected
