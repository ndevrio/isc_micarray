-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
X1Zkh3PYBPJPH91JCz9BbpYI/d8u0gROO2403jJ7MimvXKKwZWWB7dnFiuJjtGuG
rDE09A3lVYrEHHOQ3YTtbBo1esw329tVQR+t1Cas8eddqErzDDXBQt5uE/Bif6XL
w9yLYAneJ6enOS1LWVyc9Tpqvm6BA+l0p1LwwJJaOu8=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 7785)

`protect DATA_BLOCK
jCWrT7A77y9uj2y6vtRFP4IHzuKn2VAGe48/cUy670gUKD0X+VzK3wfznnZyckXN
TR3KjCNktHXGdpVfz/vNkSi3f7+TGcjGYsgAmRWKt1vaCyzkiYQeBBpwh1qToS9D
5ROzmKDfzK9sbz3eP1IBuvbQ0WKnTsOD4Q6vEUXa7Q1Q6XU93wxW7EauQlkxqOiO
csLzmy1YdsFo4/caa0RNf2CGPFBxw5helwvNT3s0lb0w+eCyT5N3HutMkvZEXuhy
YzP8a+shWh9BiPm4Bv3o5qGgR7lLAi/zoAnI2QYxTLARKhTSmKBGwWbRgyMHMF1Q
m31U8gGxRaxsAQhEmqDTaRBUtz4YGe/275b15JslHRN6AiiDxJPl0aah1VZ7blo/
SEcJFIrn2jjwKsDpR8QnkZwbbjswVHz1x4cUkCb1r8uQk0IAuo9ZVzzIP+pDz6dE
J7dxTzKVmu8QWS4KBFyNIa3MC0xU+7gR3O6M8UeSDB+MEt969z6RhucDrUyM9bh0
kP+0Ako75n4dG1vJzFJvvUeBO3ncnRmpm0hbI+kg6OI+xWyWF4bbZ5KgvunrYkAn
1bvfSzbV7m5JPytocCsec8oLzhBBfsuUEdZEfQWQIesVLt9fhNoZ0cfKz8uq64y1
tcfNRqkcaHx1YOz0JoZFbad9Fa/LgfjL1B/awBQRExliauQpT2kWlK6xORVGsrSb
Uiq/rZ9GGlzlnDCxHrJJ5Hbq6xGXBboDICnlBtymyWSHfI9JviGumE40AjbHZja1
ZW9J0H8CJQ86rCdBYEwWk9kIBnYaJiAScZBZZ0GqppD6wysR3fAAzYyItqBpIE14
Z3CqgBHebVM5Yk1atkFDrmvjrh+3fpvccNILWZ5x4i5foaHC752OHeBXcxjvSPn7
6pQycX+zxrK3SfEG5jiPwqjHoH1n/Nwg2k4RERGPlytmJUye54bt5t+MdpVzRucO
8pH7xHKXXc0iCHnKDXbnP77XVMn6aCvkTLlac304wpg8EkPpZRftWhNzSkxzKAOT
uIE5763x2acMBKztuyGFHptfr26o/s3mq2tBDLkOhhJhARNtz06JZHk9r73tmIBX
dwKSQPhL4BmEE82y32BPixszBQMCOPR5wjTlljoNGHJ3Tcc+RO5Q+1DZBVDPxR4F
SF1uQCzbdRh53CFRfFjteGGBos1UQSwWNaJK2WnRuBS2XHjpGKAaN5TJNWoEoUEe
HGSukFUGvGJBEYHBFpnaYdaTnldFAoRwkKgXV1vBrO7I0P9Eha350ZbpHJHuPfMC
QDlW7W5TIP/xOBRPJ1rezEquezOmmfEahupxzG/Inj2d0mzE7KmLNitLIhwurJ1O
zYtvhEspwbwuzSgaJ1Jgd8BJDaXUrcMK54jseuaT44hOxLaNQd840cxH7he7v/bb
Qigd3rc3qAvqCo2+kG+NW4/UOihMnRbWkMVX+khvhRD1ub+qMGJzwpCPoaQXkmR6
FXimH+PhSrNDZCMzjuihEsZk6UA9cBnaxuIDjz+vNlUAzPyqQIzy5c+NSdL2gGAf
SBFLXUEwjVQ2Na7W4DOesNMtqsLab9RDHOKen3ARlEAZflqZnCz63d+T0BzfCqKe
fU4srfViVjSZXc8JJEzFCvIS7vr8ksEHaazOo67ZJlU9TwlQQKLoTixDQ3XMEBmG
5hpLUJENugDnTGWmezVWB2nEIjpvR75OTR/9mz8VxAByo7da16Wl00RZXRsNKTcp
uL3YNq0UrCbBvVGAK1R4gYhGvf2KhsRBNybAGiWnc0wCgr7bcNRZztlqb6W4sq5n
8cVony2yDXRuF/YHDhqHpy8g6avQ+ei8owoJBfv1vUvjSxCbvw6tK0ETA085no4E
2gWoZAXmapdph+n6gWNf4db2iC90k0NRR9HBECJpwSMD0YFvxXPGQOecGgzZEXGx
e8onY3FgnrsewWkYBjvh6DyHfRfOKIfibG5G6/Is2ZZbmemQTG8UkEBvwb7DmxXp
kDdRLld3+J7PGIjRQo+mB6P5AdVd5bxwqmvePqcuu3Up+khnEX/pIVQf1jXiY0en
+lP9DfYswJXWMpuQeMAXyLpR5Xf1vVuVzzm88Po55TtqcPcyHkn08M5BymZxNYBv
jKhukFxcdbL8h+WrCTIRsF6Y9VkNeFLpZD73P0xa/HCrL2vCitB/7BFodwHzLX7E
joagWL4fxljsuMRbbNN1qyEDKqHpdeJlAsUX4NSSU9S4QKkl1ugPEDI6ZzO//pDA
2UnPXHFhPrLiBXzPSvalFKDkAhGdnL98iN7odhdghHSfaoCC8JcBD2+CXG2ajS8d
pzCo6STBjOOFISt2o8tBEViAwWrl9CQ/eeqp5pQaLnwYcHJMOPGxt2it6WlrqA4M
CBaYsPQpX5VnOO/c+PyZJ3mXiuKjRJVOaj23n81pqDlnBj3sjvXNQHx5LNXORVJF
+veK0BYim++wCzTRtAsQvmNNvjyvIV35k0/b0Qxe53RC4UUVZEfYGKPCdp63uMEJ
awI1CbmrvKI4moriyfGCizdOijiKL9Ni85mMiJQQKiGc0o1FZDhXOaKMvtaVNRxV
4vU7ac660w0/+uYs8LbD/nBmiKLr5GLq9gZE7EG5d+YcA42wztP/fFf1lchoi+Lc
3VdFvMgy/fZupsFcAkbLmwfWKmCfATjR2fb/GNg/vALGc0Zv+4tKR4qzES3c10d5
wYKvXtA4N5RNSx/pldwup6q9Q4ZYRyCO5LBqhe14cyLukU3jnU0KmTTRw3Cwqhzk
NqPCuyViBj5vxnmr3N0Dd3M0m9i6NXmBnnL9aMhTLI2PUfxwh8BfpzC+Ih5TGZEW
KVqTch2FnWkf26cgiiwq1hYhvRlbsvSLe/QeAQOJOxFfr6jyNR1cSftIjSMJlkeD
wvQ4aMjvslQDmYTB4sI3wXWHGGl0rvjDPPu18Xivz0Q3NRRKWtp6ryInnQE/HCaX
fdSdSjc3+dCwCxH6l5A+IYFahCw7/WkDXZPRACiflLHKkC2cVkGhyYjVDaoO50or
sGRZ4EBBpDaku3psUu9iuTT1zOdUsAVNjyrVncWZT7Juugt8/9LoUrvMP1JFvzVJ
E+fvVy7UnerKXErQQ9En6AiOgcuZZbK4CkHt7CT17ArCUKTjRjrqFLtb4nWBph4N
cjF61pkHdYVvg8w5SdeV2NWRWLj/2eKWqV4Nkaa7aDSiYVIa9sQRjkmNqemI8nIq
i9LRiwzbMh+YX20USYj1MX1J5NLw4PciigXPrPO+bAIiZdk5R3myuEWC7pEE1dC3
GKKDlDUdCdrSJ7aZA+ngVQQ1hvzWbGtuXUUPTTdiFo7pt1idi2KX8Vayjhy7QmF+
ROGjcXvdtL2T2H+TmIzHTv25ClVDm8c9x5flRfekQNlx9D9kyC7zNNcG6zHZ/crW
gvnp62EUbq59PFSqChPA7j6fzJnp1nk1MbN+tYabIJm7frOql6GfyAPkr7DF5jYn
2Dfb2axzGMAWOdTdKfdtMa7weUJDh03N2SAJMw+ANxQuzb37eeqpH4sIwlWy3I8D
se8+hjxKsudS63HfuJvK2/USqSFUf9SFAbL+ievuONKWslsUk1EQCxHCoQMVn9r3
hRyH8GN2Jdi3HI4rkjp1rB7aRQC/5unbeGa90bJUqGN3aRj9glvdd00cXpEEMH6K
rHudAzqJUUn2Mg4/3A2HKxHkSC8Srjr52vvmTUSlyubksN0I83BzUAv5K+QDnbE4
DrCWZhmsKD/qXPc2xqTNkPzux6l2t72PS+I4sOlGmsx+iZAvM/pJ1eWegz83N84X
MTFGAUwxVd3Pi4lOG0TSCv0Zbc6GcSl8+/xvKc7jjBL5qmSE3ePWkiguxyG7X3bM
iilv3Byf0hmgF9G0oX7oztlHyOnOIduDmA3C7T5ZuP5HnVrXOeySHbrRCbTNfglY
UPbQQeXE1CKQMFaky55YIvsYHgCPOYYWOzRnQSDjldZraQaaeueHeIkM2wYIAL2O
ZAlm9uZfqZUrnyDEsLsbMhLx0VS3KTmAiow2uojiTcs5Wo9ihUJPqUdFs2qX6XCe
3lN255pXT1UXdA337awJrdzyomjAP1LeTa3Lc+9v5qqNvfpreLH9kmqzms4Qf/0s
YKrKY7rkHqq1fyQWmh3EN+Z26JzkHW2Eo/0qSsdRulyILvlFin9jwV2vHOiF5xd1
mIoT2kcGa/fT9lMAFQw75xjtDpvrYuto0/W3/31NISFYCzyX7SNqOK0TIr6so34b
cSC55gIkmm6iSC54UXSSOwIbaDpbL0PKq81BjkWZeDf75WvTbcs/UzlxGL5N2ZuY
qSiQEL8/o+z8+AZlW7Lj9XJ9oBeqjSRCi6iMvqWTmIb6xK4r1AXHaro9nEWwxY+A
QbM79uZpHW8EyFaiv7qvW6sAg1ZvAkU3eJFEftLniczQl9v3DpL8a/21tayEnwlV
G0U9SWoxMyHa8EUs6tnQSJxK3/6p57rIer45kJnhFrQh8PLDogVjmbpWStQiX4P5
8ztjuAa6/LeY9znB1sdVw3pKwaU1JV2ucwMyrtfe7ovwTAtNrJyt//7wvSKEy8hu
UM0obZENTLcUVilrUDONIVJEIms0dwh9COS8Hkml4u5wtSX2E3WnizFsobfKov2l
I+LNufuuYEZnqeW1zdu9aqiNRNQgi+Vmh4J4Mzg4e39ggkKWfIUNJdHav4VEMsdh
LHZk678ss5CC2N53810Eef1BD+WBf/i4s5H0iX1zzdBsp7oxlyIi+e5hfgPorg/e
r2cNKFAjm2wieKSz20O5BC5zQcbPRTj61nhDAnhQmFdvcSj7QprLERgWRpx2HOE2
KBJD8uYqwoxZYdqZT6O5FVePA3sAKLtJnY0aUP7K+Nsxy9VhH2RacSA45o7PflA+
jtGgQDIAHRWYc4uNH4TlHuz2N5H22mQguI5gm8GNHPwmDNR4NzCuRiE/LzyxBHlU
r5xZ7g/ey9wi7j2uHAnpSh6ZoZu7U3QRdeHBg8ebRBztlyxLK2EZDwbUwQ1UgzGx
oYcLK9MetXpglV9RQq1gvo2Qh4r05gNtNqX4CNv3SVRaTLLS8jFUVPyaL7HOnrmc
t+QZrI2oXYdtV3qHLehoGemB0jMvxco7vajqFsyL7AhANsy16ocA3Biq3Y8KTx8k
XK50zZmKe4SkZEbGwP1Vt5ywyIn7u0xQLo6dqYj0jRxBZHUPrtDg173XUE1+OmCE
aST3NKteV15XNf6qFB8MlKjPR/LZn1/t5I8PVZGBQ44S0gCfa+7mjqO65bD03owE
bJQRo2kZq7VoJb04fQKRFianDJ9ot6xOMqELYe033kLJcsCLsjFkyqqxu8sblxwr
VmtFUh5k16IRkqjdT8mCUwI+OD59xaYgumDWjlteGZ/dsq/yHPEo3/2jAqHbhN2I
yxTE4klE4Cy9E37KGDKfFifvUT8V/Ck83ZN2uuq9vBW6QosmYxMoXYh3f40i4Ia/
g1R1S8x6IetF4KKOgijgXjC9w1tIbk151jLWhV/GjFq/2AyxlnDkNxFwKdOf3G64
tCZZiQF5PT7eYT7rz6ORcXOuskHEJoSJO9AF5Va1MPIkqRhblJew/C6M0bbBa+QL
//NagX9EsTysnWyDlQ4wk5VNcK9B+zzvyXjWMkQHwOCr5jBTt5ryJdRWW24LU+3E
vRiaVwG3Z67hrYLQNO1ZmPPo+h9EG+yrH1pfm5c74WY1QpNk6JiN0hsFEeGlbl4y
30xH97Kyu9VCwKVCmmXbdSDtPtRpGiqmFqvKpMKdxU8aVb+0zUJ8ils8BaOP18gM
X14YfXZc3wfhGdODmVjAI8J/2GyHP1vbqOYYF/JtRyxOBhwzmHJdS18b4lzA4CVX
uhL5jv6qYk24g9YLVi8cgBSLUopfbeSEw/kZYRC5WeL4TZZlLjk591FJRQanjLB4
IhGWVWJiUqjP6mDtEfHYeLqzWHFuiQDYuVr73xdyHH0GZwrYfglY++EftmtlHLMz
0fX6UG7ezuLFX/XmDRsLkNcdqmR1lOTIU76wgQGemuoK0MhL6WmPnzuHPtto3/Lm
iYRi2WyvCfmBWlWruXqDkPHQX26trEAuXnG0qAnpbFNFHg42rWt+ldf2j+WW7EOw
oScUpPlsLZLrXf3cLa8Ar4EWPM0efiR5kO8jh9BErB2NP5kX+2RP74mhBPo9NKRI
yS2Lw8DTPUFf1fdazj5/RtZFjHGm3w39zGGfBt1EF+StV+YII4/leFEqD6Z4qHep
QxRdQ2Md26WjM9gkmTZnb9lXECe3LfsthmSSMTjsPvH3O6qUPjOxP1MSOsto46DY
dfADC6vS6ftSvAnEMD0xLjehmJPNp8aVMc8KrE/xcipcZjJEj7BhHvZbn59iT+uv
h9x743vtsabigS+UQI2MuP6FtrKnH1H+xlPwBlxo339B3WXpsswGsmqN8rfXxovp
UBBLjTgZAGzDv6hkOBqP/MSBahSmPb5v3D/vB476YiH+lbLZgD/UVXTA1slFvZK7
1VNIGHhGJTNz2I+KNqkkvQGM0LEEcIykBg8J+SZGVjqo2HuXQ1BHcQsjwAPUT42G
fiMmkYsOwM86KLCAF3WKp3zdIpE7lPDhyHC+ReSnVpeFKBkMaapo3wk2ROcVpIuk
Brpezu4kypFTYmT2W0GcxYrBZb2/5eqwD3VKTlR7xDoSrYGrzbTiVR6O1neF1X8L
WDd0THJtCzRxdXi2fAgg4LvBBb9ngQBOJBpm1ujXx3jtM6n/sIujxP0pymM0XLmv
JnmmxsM4cq0sg7SOjn3hKFYgZmReYo/Y43R7mZQMqJCHVz3M8QYJyTTzT4NL4oqH
NdG+6u03F89zCn0g3MCCkqW9we/73Vzc2jzVE/Yojz/dQceG80iqmIoH4RT9rf3I
PabcweMYtKiFX+BEWi1PCtBQDYShQIxBTmbEbIDVqSAPoJwnC34ZPGJ7Tk3OdVdq
bP71i9bgYq30bjJZlDFakAxtLndmkIlBafFVzWXxT9/FgnAVj9ey5DWfE+HZ+fgO
zPrEM537IqgSI7fNo+Zh1bf/hjF3Zl7mOZfXe3UUC9QGSko3eOvFEmA8bmj/lluv
QFdszmpygmVCTijeWNg7lUWbwBHNW/hbJ72bDR3diXWz9Wmn/U+kE9FumIJLALos
9J81KRR9AQfXLaKSJzVeFlqv8rEY+UTJIDTR2onwMDdFAmnaIHW3NOrFGwW8ud46
GePdKuND4ADcM8OlZuOg2AaWukBt70nZkje2vZTdcwdpwBuJ+W/8sHjTSqMn1zNv
mx4ZCjSNM54BAP9S9pWxOrdjLEuD3h4SGdRu9PxGOF50WRyTNL65lldWbpQ/OifG
RBI7j5GnsxjkZ8smq1ZZSqfU//nVkTcw2wp9ovyKMV4IDYPFY4rFI0nCxl106V7Z
SQwmY0gZMohER7gAKou5K8I+WGAsQz9pn5hviCH+ahPA/HEAoN1Kkde7S4IMdCKR
rYLbHH7DWpOv3ogyPOnRE7Gbqi214MxYDZE1dmd3vDaCcDxF4Xy3QkIvvX86wRte
QNAyxvIXSf7Fcs+VL2J47Hiq+HHtn9s9jhhd8/SdzNdeANLpX6DafIIJ4OAvm6g6
JlhHC0/zjJnxCa9yqNrsS6doIcvck0ZMEZ6F3UBOZUoM7QUipI2Ba2qW6vEUrkhH
14WG55t5+f52zvp7AMJXYjhmqPSEQV64zOEq0N35Gt0nbBJORSEMnNJ1gcse8LcE
QnuvESQyTunWZUIuspeQ+BY4gACQf7aRVPmMdfFjvMqQ6BZEw5ngX2RtdHhJPsW0
ti36Sh9qrj/AWiQn0HvlLhO7iv4+/mexfoxgLipWl+R8oztdEDUX6kG0ygp+T6LW
9dZu77Xr0x0MpC2AcESVcphkG6Ag2XYVl1NjsCYuA93n3UC4aFWcgMXI9I9YmoGK
wg9Wx2jh05z1ICobGXCtHGOPYtkmUEwkwYla7a/f8hoczz1Y9NRK/867qUeOf98P
R4C5unMJLjZ6RZRzbCBwdZIgu/mhhYZhPvw099sYfYE3RgqMyWneJu6Xh+Zdkwqr
43dJyywBhfpCjGCEvnfh4G5sdMZjJhpxLB392iMRHQ0xJY785/3qgCtiBKtCqy7J
loqy6SlZQNKKwzwSxOOzWTrNxRasQ7Lubc2b0ZagQXuk//3DwBJbh+noK45DicFN
1kWIYZDVVQV4bSrq52Mnn1Q0414oRrdmMPxrCbNTt/eVPVTDQY4576heOAM4BmaE
8/zYt8zbczQ3NZueowVlTjbnpSlgRQmhR4yGHwkPmvbmcy+jgPQVIDMjzw8eCrcS
j0+aaJMDqWay/uthTbt+tqVpOIaFkuyRR2uPZOrZF7EFj4b6kxEhRYz+sowJS/qW
iezN0eINZ3UwB6seTrcL5J3fPdMEAowKhzekKnhad+MKi1tmxz3q2PHbp5Ve67DC
fP+axP60LWRtdbFEX/XMhI5WknhKbTsiFtj2Kfqoeyogn0H1gN5m7cV4IFifBmTM
S8AGYzQCsGGM3vwFW/w7vaIjJE5Vng5TQXtiiJhOKFy4YVnZ673lT2lBQb1GfBBD
l/Mx6joUR8bOcZ6yWCYvUhZBE65wBSrox0e4QO7MJGXu67a4JrXO1+4CwtflT/UM
eHsuPa+MSFl3i5HmEldaHw/urjr0D8m3dF1G79QT0dimBULrfWLL8akbcPwUKf4D
4aF8WHVKwug+7BnQY9OkrXuN+GyWHGRms56GKX3tLr9yTY7a3TcukdOdhLuciFTJ
X9fAe1PC3OXZdcNrtHu2Ujw+MQtYOuO99+OvL3V3jpeNamxjmlTYYaU+OhYOxewv
aG3EqeFZN+rYiU0so6nqTSitobeS+tNj4TVqlN7epDWPRK2P2D8kyWYsUVPAdsXQ
VCJMYU2EqMBGnmSodkcs2HAEVuk0ljcu5nlOgTsIYaPqgf+A5iG/OSt/oZoAanFl
X1sY+/vHvpUBMcSVoYsihJvDaD5KEXRimGVrwz11oOSdz069faBHNpVlFdc+Q7pB
42007G5Re/zGKtq3n40tZ5am6IfUuDhMl5GiEnDyYDxzSOUmAeshgV55BrgiZOIM
FqaW7rYpYBP2Z/ruAPhNCtzaBkTvbcDa3zpQNbNrE35QBAR4TccEBBouWp3CjYe3
nEYNzJOfIHb5Bv4X3Ja3sko279dEMmsg3rKLlzy4vq/s3G7J5xJbnjdNh55cMu9W
eu6g/fshbraxjmn4Xzp6m/76pjw2P0D/rOy3jTJHXeBlFEtIUMaTivlk2zQkZz0o
CcSl7UWMG8Cq2EcpsWagy1v42chL3y3YeTbcMO+wqQ2NnK1/kBJVSWz7Bfu5ldAi
V5sQ8690S0rdigTt2Tf3YdopvUt1/iABhCTGdrSeOwZVTIHuwLv0tmig5wMEblTC
gXXlOFyiDMADgwBW73UJPjAMpyAFE9BHqVz+Y2ozCs9tdyQsYf5AvsjsaOyN/O+c
6iqezjT4BuU/USnGbqD/LVcXmi/4IbPnNY4i/3MnSIei1TP454i8Rqhrv5RnKAwQ
Ywef72fQNsQOA94Uc27siY5Kikv5GsdEDmZ3/MH6nTapGHPN+Et3bUpQWBbGX2vx
Xk7nFKh+UYL3jB0m38/VmcE7NirkWfaSuIqER9oso9ZTB2yxZVDsm2+W5APy2S/4
67tZIEPqrkSaOb38a0woG8Cr/OA6HgkAJQ9B+Lv5yQ3i7PbG2DlpjxiGnFEtQ2zk
AvcUS8bQUPVXMYsdR0d8KcfCLhL2GeL1Zd3fWRZpTaBFfxTWGayu16zvuMBRyJs/
/VjWYQDP4UVNBnhI4yDSGdZQtygNRKETAeVlSAxC7tozXSTrjb3QoEUGzKjszzmj
ARfXCGfWhxosfHENimyfSff+V0uUR6cO0HnCNnHHFehjmBS70QO42X5TZjasVhNj
feqJJkIL+X0YLXFr+MFtQpi6u/OiPS1PFZrqMt8LG9R7cckrO8ktPqLRqZT10V1a
37bYAAcBZzyS4WDJH025Xd4EdMfu60FM2RDp/xVCuQXh398k6wThVY/ygapS5j6O
4Pcx3/i9Gy//lxdI5Q1tkhveAq//QDE69WJoAilP3wkTcq8juG3LMqtgF1EdKPON
xNtAGDZbJloylAJFunzJb+cR8zyBKfmqyLdEux0EDFOB3YzAVzb4QkoDztLByOa1
GtOOk/BwSjE3e2rdr9JqzaoWQk3NQ0pStGjVvaJ7R6a+5/qyKA/A42n5sqkEKLA1
2IMiVKaedwwLwnel1+GJfKlD4ufNNqtn8nX97DPhtcE30Yg2H6tlR61znMq3g3bb
tcC5g/owq+QoyPT2CTFYWRePmc6hrH8VEEK2qe8q2d0B7J5lJpC9Sk0t232YxJng
DyAtkfdafzn9ubfLys3MPNaqonbU70QBW4zAJPy9okbSvfB0XXc2ujJa6Z0G82Gt
hLGkYUI4QMAKprUSrPRp6gE/52d7IvKegirU5h/Z/4A=
`protect END_PROTECTED