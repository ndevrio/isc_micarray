-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
UD9xuyj31TLcb7Mlk0cyzR6AROado/48eDF8iid8rZKNCNeLDwIiIrTJ6wxFIg3Q
JX4QeiK/oa5JVX16YOzKcx5RHDrdXiN00ItqfkLo9V1+5DGwFGG5J9hSKbaNN+Qc
hdJgMEGe4qIPN1mG/hvSnDl5IbMI4G/7d1yygfdIqlA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 6479)

`protect DATA_BLOCK
HVKn6L9nNw4rnDUIAiGljy7rJse7fxxFxMNK00tUObXwhK42W6ZsAQpfl+Kv63MZ
qawlNYGbBoKYgPjd+Mv/zBDUeLd5CVKZuydoPvy2px3tfJpPX8WZyvFmYcbjs+yj
Vmc2Y3yyJIBSzzxFXTPFxbC/vZM13+w7UC2Cotxq0Re68KKey8NRMQh5A5Eubdil
NzkOdR5tG8pAzrlmpv+uDVkfl4a5CO2tZqQX4jUiQgdlRuYYykUVBtqYVuqxoZzM
746QU3LAHakcqXB8UuVwrHud3Qf567SsuorI+hq+fRFfKtUmKiqbQAZFc+b3UaZr
5v75FiQhOLzvzIxPfhXyy9xArnUotaddVORrR4iV696bzuqiXEAxJL6FjIeSzCYQ
obEIgE1rnFf8mx6dnBFi45z0ATYI+PgkWrisRiI1VFk2ZaUx+IU1djfHhjw6XU4U
40iyqy69cTN0XEpc2XFpYif7J/F1OIcQ0WCsyj9g4EBqIwyD7ISdGiOw1hp1XphQ
xQgtlKpj5bV2uul5DnZ5QV4X593i+1BinViXP22om07kWrXcBwriej/C17mMyxy/
SM8FuFdNVkt+MS6z1qPwGVF9UmQje5i7KilbKeITyJPPokEYFpNpBT6Bx+BrD6An
OZruL9hB53181kx136SFW+4+HuCtgFw7Lsbj5n+8y4UwEJ9sqm1UQO8r9+mfgIQ7
qHY+EuBHQa6bm1aaS77tVD92LKSa4+L6BCu7uyxJucyBp0Ze1O4dun19TbK7j5XM
l/9+YaNnrDs/TAuveITYwziXrwFoduxvkA8oUWToKWCNm5mJfl2j25NXaVXr0bP3
xGCZtRChIH/Qi0PmGTU4S3tz7Yckms4ryEZnfvM2/1S9osvD1MVfsn5jT56OY6iP
LSiJeaHuuEamdN/UdGCX1UfXZlPXbRFt1iLvA53kEanymK0xU8UbXgGWsTSIZRP6
J48ptLe3LDwRj08XCMaUAxPLcyWpJKs7LtAgW40QRZtRpwgGqoBhisGCOY95q/+Y
ajfz4l0yH+qcc7rSpNGjPwfeohz+klQmKgiP2muemxPGqYeOKKYGuFsYbHfezvm+
62fMugp7WkyhCeiB7UmKTKNzFYhYjpi0cIcV/CDLn4YdrsJNBF3k0FbeGjE27pTF
MO3V/6veCmIPdTv/ydOiFVYtdDVxLAcSouZRzDD0OMMZdUnQ0ALnYo6I2fXnvnfl
8cTUPx0VjiTiK5VHNkpdpgbLzw5Py2szfHO8WyJqrd6aXZlLZvpyqDQrht3XRbm8
C5HMxDZvOF7ZJ5FPakLQnQNRJBolB/mJvppIRfUX7LnbxGrl4mfUsbwOn5vmomkn
7a4w66o1KNRh866C7DQQ2aYhHdMbVmBDgCIc7j/apAYl0Nsv1umpcWxFCQE5QSE/
AGu49PRvfnAq/Wwo687JaVthhnknerCPgcI/gjyXhbMm3SWvn0NEziAnsefCSQ0H
vZIiSavC1jDxF4XiLMD51xq9X78k9S8GkrQRnD5VP7F1wjNz+1IXZ9Xngh6Vo82H
fgEGpKS57LmBuVJDgFIFiuDbbBZIJGUDWFS0CYRhNlANT6SCS7cdjM3VM1twE3Nz
CeF5L6CX7babIi3m+CTHl8pdKDEprcSvzkTkU8i47JrLvJQJhMmJSjLMe8j0MkeI
A52nTAOk9jjRAum0rmDEyy1OSC8nj5SrXZCU81+jDqKofk9WafOS4a7RTJW/osqj
L8HprhFXAl1OLhf9jrEJmpABCygaApmeyhXC6aPjoEaN1w75KXsJbqp97/fiI/bP
vwY6NEHXaHdNVlM5Gnvrl2YgNSCxTGKSrRMVAbI/J6HFIcP0UuVBrlxWAMboLV1O
GXLRj0QeLqpM3ByWmwGc4UKxnRPrkJ9oDOIE1J0AKQXcanmaiMaG+lXcbpz9MLqD
1No0sVdDm/PXkNGItGvJSvV/UJF9arabbXslI3jnVCwpanQJLDIhSlEZFIhR0AGL
XPIk56HssrxbJKqrUuwLvG3VuiW5K3TYe8VBiiG3wn0XPZ6f6qgGjaoui+CdTXYW
EOU3qJcDC1bKRIT7xMxiGezVkhE6euRHX2cnKzIHoSMs/5om2DwS0Cct6EJ+EpZz
kgFHU+VvcK9TTiMuUWQcbfngfyK8pSyAlXGWy+6xXcdptBKV3uPY1lIdMnEt+mDl
O1L5fRZ147TLI3B5xc7qr8S8gQd21zLr1L4k0a76hKRoSyw9i29nJ0eozEtg01r0
CKJZLML9USmEEwPeoSeA5I3Id2tkkL8aHK/yhtnDynbswbgkR5YADdSHREMRRs5S
pCUasCSVwN8Dkjpv72if+v6AsgF3av9MrogN72I5n97u10mEF/C1vubkrQlrblAX
UyjxJp9p16ZWxGH/aAA8dlP1M+BJSnmBoYjfpSIwNZ4bR6SZsmcJ2TLfUhYuSTFv
xH3AETzoEpu41V9ftWm4vEDKO6b3S0dhiFSMfpynyefFUXgPmZAXpZnShC0HkCj9
g9R8B91ZHeXYTELa9yhz4gYLOkl1Oe7EM9I9WBBcjbYJX/LqKAfiniw8rAci5kZ/
Tb4WXXFK3HVQCydi5WByg/zxnPpBwtuX49/ETL2v3NMAj0mdrdutefBsV3b3nN4I
Bq+yqLu5gXuWmCSwki3VBKNcFpYhF8CTqjoDRnu7QoH2Mh0FsKhoaatriB43YYEU
U1SkcPfAYOXL5sNfrnYQ4+S7JoY+UHI82f9/VuCuzuc5yhbKdC1kiLtnLPwEGMAy
zB6OuEOJkqggGDyZk7OH5kA64DwdLN4oBI4E0X3hTEKfaIva6yN3+aJDfCE5qLEK
KrktEeWIfUNNF1ijENqIviWEh49ueD5OXMhDYtBWHzzy6rbWuTPSvH9wD+ZlXiyP
fmNypLEKGtKbPpJT8X1FPOuvaG9gDvLg+ffTzGb7RgBl/2evkztsXK6ulvankXe/
LDEwV8TjM9hSB4pE7cgAXA34NKpByScUZdhpkCRDng+H7ye6ARLPEhBCIdIMvMEV
leC+MG68hYAEkEP2SDK6cKZFhkQWmm0anczDll7Dl/iO8MDH8YNYNoMmQieYc3Bt
Oz+uLL7cJncF9mbXIabgOm5kkf+AcHjknRsfRPEo1aPbG0SOh/1skm9etMTWi33N
TpZBvBAy5x1/Yy83JwYTGSIdwpll1X/qjQC9xzHl1V7UEFMfoUQNF8J0DQRH8iUU
DFVVFF5ox9twTGtSZOI5zwCnDVkRDtQ9XOg0OGRKOqxze5WUeHgZU0m0QWps+J5O
mz7iNo3rcIrl0kdNqUOk6BEDjWkIxQYTVfqYMIZamoFikJajBRSpheRKoj9M/6kF
0rNzLF3MsSZRodn3iSHvG7toVUsakeciOoEf80gbTW6KynPO056M6r5pjfwAisJa
BPz6ptgggylMLX6SqYo8v/yt//xJtHkvHE7OoukpGJkg4A40sC5VwGazybfNGU/h
GcSm2v0/lKJ4Qskz23AG8i2R2Mo+eAv0fuJW52kuE0feWgj+zG4Ngd9hKhofteXn
mPVrz6zmEY3DyHP/QtHP6Cue4UenHrqWOdJ70k49hm1Ae/Olx4DXiNM/a6KGJIhb
6Twvi+iGTsQ/I0t2jXjMbv1J/66v0pfO5HBp4iijaFs6P3aEhC6NaH4+qHpzAX3g
y32WagI8M0mPvAVburUtpmDApRt1SvqBpfVwl4pCY3hqu/N4Ta6pl9rfBApgZ+LG
ZIlRx2bRvJAwZvl0nQQFJrNo7LYZ/o5XhPM/mlN1RS7cUcTi1rCsgwYKdqEPMvNe
Jw3DXOvtdBZ0doYVMG5EDphrwa1zgqWhqRPstgN1SCLLK3vu0uOr56BI6CDIRyoK
NO7GXNx3/0K48fSJCZoJHT3mu2A59m+Bnx9VtjuiWEoR0/64Em0Fa7SB9TysugaM
XUp5v9UCmmHcOY3hDhIcRpYAHxJqGLYvrRg/xzP5X3BfWhwZ/fHSdWYN3fKKh0ic
mdKtteecvW9iNm03qFI1Vug5ducGKH8EgYBxW5+aIwpoQj+BtLo9YH+WT0x1wcll
jAWPf6nJ7siY7yiLjMKL46ldst6qZByLWy2jb/ivkI5pi91Gpn4L0fC1byDTL5Ca
t3gdETARMufCI548xC7nE6LLRuOc4IChrN26GAaLrdWKXNXcAjvV8RXJdACmRm0N
ztY4ON1f37HrylEcmxEqSVYbOm7M5yZ7H5nC+xPH8VfH04e04szsLibIVGimyD1V
eX3E6z/6jebLUfqHbjNNgae90NjnQocHbxrvzo54S+f1XCYuc19vRV5YWp7McWhn
2DU7FTZfnTC05m5zXjg4OtG+hvOnUyQhgIhTcp0O8nDoIMxaXQDT+5YFWl7eHNq5
zpy7eGqtyoBzqkiqkMlP4tZ840PEbbaK9nQtpUqJ+k1tx2ejCEeO+lgF64DBL4GT
5hbb7bxCSBAu9Q9wr1VlJbXqNuuOW8PlBIj2uvxqPCJHLYjnnPf7JSAiTY06nMZP
gnlUYtcVTGQl89F1Z3OSQReJ/7zoniwbo9AmM/hnw3QW72YPHgBEybX6He/2vOI5
F2BFs+VYGFLxl2oQY1PtVdy250a49KmLBYGglCBB1XE3FF1pO2owYICzFJ2yLHah
lpfQMq0p05DI7qQVGVvW9rqPJGGRizH5/9QMsyIF41PAkCvpj5NqTZDI5SfYUgzk
4QfGpMFuI4YI7Tvb9QHokrZ3fNSHCiFz0PMpZdPnV+/HO/Ddsh3kiWoi028pwYsv
gxGhfMLdexIx7hU6ib6kv8Jx2Axb26GoBz9TREa6FdhgoxLkQcncHA8/h/Uu/rB6
UYHNWSURHduihOhOJG7PI05oLHwfnSZya1F4D6DMXDkfom70ruHLQ3kXqPmU8bOT
mU8aIsy9fxI/WgDyQ93hhHeruSnpCrS9r+zyol61mHXQ6tBqiqrwDAK1NgWdjW3U
AweI9HBKhy6yeySYb0th59E3ka0nz8OCvA3q2UED9CX9GayIStWL661qAYND83QZ
r0eMqNrLzB2yVvVtuwT1uo3qGaIOEzEHz9Syqnt+m+Rh4TtfnVt0tpH+IAYwAyWl
K8L8BFJY1s7Aqj6k9qJuCawPZuhb1OFn1yq7wL6CVG66gWBplqiwaSf2G1T1oc4P
NZ7YhYVb4V7HRCgfo2MedYrXOZ8gCaW/hEifNlgj2U4yAcUQluhXuqhIev1RjyOR
OI7GRub5dgEBjDNcrG7W8GNB68in8/jaUwVuiaMO7oqNpt9SGyIk8u6z6TYfQ6mv
uCXGZwXdAT56ecFdgipyXBuRlwxre7Kpf+b9Q1ffLN0E2zHwaAjk1Y6hbGuqDcs/
uFl8YgjfmPbpAt7K/uxblaNIm+do6gGjqDzELpPmpb9+XiBbAVTjAB787JdRsuVu
h+fV/1v2GWJW730GzYWbJGgRKnSohS5Gtxt7JmGwt0xvx2PWhZx8QsiboZvny/bL
D6WcoFkEV9/abLcVYqcemelZ/UkzHY5W+p7+0WHekz1JeswhsDg0ZuonhENLvzln
FCYHx+ABbeu8XYbIewfhyvb1lKYQ8Pr4vJayRikZqbyVrg1pcxAOfsZQiZPdZTq5
MkvPZAAS+8Koeug/gjdkH7oP8vqbsurVG6WzVsohhCN2hJA9XHRYvxM9yuTf+HEi
ukS+GMykp2gaanjkXeKk5VDphzhvgKiU1tiJHwjglybvGuZpZOAWg+WyzpQNs1ic
PmT29o6SMjN3H+J4fdW8oYD6Y26c5omlF48WbL8IRtOaPS7Yo1jcQoXzj85N1VuZ
12lZTKUZ8xMm3PVVInnAjjtViNFmDHapGv8TTYahdZ7acueiIumKeDyl9DQ9ZCOM
80eHBbmBOGmivG7NaX09VCv98QSJDYDbx5FP820exEQru+AwjfR/TZ4AQEEzMWMj
fFMKdnxGzsQYgp61gGkZjEa/NfQy+Am5HP4qzlhcbUYQEgtRlHVaELIg/M+ND6xP
pLYiZHntWRU2AYs/DtHOcu/lZnh+ePKEHXrDvLDFrW4SeaF0valk8ZIbhQPcJdMm
eh44olDpkkw0dBuqXV5MxmkFts0yEgWaNPXc5dDi6OagirvLgsYgB1i9KH/sgg5Y
HKEZGmiSO6d1ak7FTJkCMNOgTyumjNQpcf1XlpojXWCIe11o08iJmAPVxkRS0SH4
z6h9sGs3ktdp8r1H+NUFlytUb74i1Q/+PO49rh3cKtCKxkvlQORWd8A8Ct+Ui1fM
+8vspYjs09C9sPzEwWzxchJ4jvO+MKlQJ6vSt51xyeIshaGcKHaPTEM8ZuGbBIlZ
1kSkLoNgfO1X2q3jMLgQoQKQlR6IjNiErKujWOK2ec/F1sVV2iG/dn2Cj2FKgZ3v
92m4b7pLuzzG3UpufO3v5Q/o1NzFefY5nS8kj3E/eZVzTQFnEIWqXNlr5KSkXFeW
Hq/JSF8eH0hydRP0YtMoTjI8MlXJcW8BoR1veV3WUsA8mub7mTkrSnmdEH7Q/BxM
WnX0uNik08nZq3PdmKPkYrCcPog4mcKuw+MXhoyVuj7Gz2+NtjwwzYNRcD7IOe8R
Us+0cDNm3IQgudCqXK9kOYK44ecXOQCFsYFUgcPyKSweqUYw8gXswtY5QUTfY5cg
B0obihEZjFWVctvVOE6BsybYj/rIdKY9TiNVc5ouM5is9/kp8DRLO4oE1B0Ed9aI
/0SG1N6OrZlAaoCjNIFqzazcdAshP6KUZ3bg81mkSGzS1+0fpRrPWkuJt2246Y6D
sTD/tOMb7DjMBmHcTKTa/v+QT+m1OiU/G8ldmZvgw6o8x+Wk0VCCRMX7EWRrXVTR
ZQyb0IOBr0ttibOEQTBGqrLWozp6AXquN8H8i290yx9RzZU0lokj7i7fzCqAXzUB
+xr9n7Hyd1YqOZ4BUkGDDKCsEz884+fjHlXbou3eu0QG0EjsfsQvWkT9V70jWIBR
563CRRRrpnjLLIVAK6VjnJX/V1Mm/aUsxNzeL7AQLNiUUPJYElrkfxQq/sef/Y4x
bKNz2dE5nrAlP9dyFyvPGzpQ/iSBsGkQj51yTMdVMUU9FpYDWQFSOu2DkJMcS7Yr
FUgxfBUUsqdchvXWft9ZMZqAGRk7bexFolH98Xi85LoFxRtRw3Q1IbDI6jWORgR+
ru4GwJP+7S/gkk9aydIIi8lCh4Glak28C3eSWqUHErfteJKkqotMGMFMM3OnLQwG
fQT9/LC8jvdvvSYRCZCvxkSHI9LuZSnDIDY9TA2jKh2q6+rSV9IaNiGH444ouGP2
NqsDNW1PQuk/SHvg+YNlcwV+B8mTIbg1tym/1KW4Lr7X7TqhY+QFu6wT1WUlqSJm
rcj69PrZLzatf9qpShSEGVJ68GB3P6utRC5L6w5UEY3nORQ5fgRCeCBkq9F3rFP+
37l5hL2CJJ4NfS1ZYN0JSSTX2YqNa4PacdbtLR7RgXcAC098s6H1FEcp8yzZQMTY
lIQLRJGwNjdETAGa6F/0yhmVvLn6y54RFpHPCA5anYv/KPctPSvvoj9bqaQIEHFp
d+FcSua90M6AhlqAp6N0Q4P3JbqXU0WYgs5z+vDZQuCf/22pEZvQAvuP3Z6bSvqY
pzyok/Fl8ZCaKKPWiUCVndHwnsBCFrJXFgDBV7Rhs+0SNoxZCM3MgXo1pgguplnE
AgRaoKiBWeo4D26lRbZarhVRBJDHUSTg5LKLGoy39cdv1YG2bBt3npKm0K2Rofnp
2yK6pYyvaXtn7jbMOuznqHrFBziEL3owsY8hzD7YTci1vgAn3aOkc81RZ4lILdKs
pa90Ror+aaCRHQld2lrUe7pgsL6krj45qt6S41I/ajyx8O6xc04UI57i/xdzhIdb
F16bTk8MeEb+AITEnMlRC2RvF7QOp+LSrLgeoepstsz2Rj8fvT43kNsSNIhxMT38
RONGT09o1pMZ5/7peMa/AOIO7/O8TNkcmHUhvXkSdZt8I3ZEDUBtM4lYFhAl5Zmy
KudkyZ6S/C25BckaxRN9ILeUvCsGUmDrNOllQ2eyU6kszKLY3CrzokfX/E8i1wpt
yQkw9qF4phg21TWAaBRkLeiIl7lVMty01x8T0fNZ4UxEjL6y6XbmhKEhmPgd3gVG
NWQFJ0EpJTmbZ9J9rlOEWm9/A7chIpX3+77lBQZdutFSdwAyKIlPlc2qDbQ/NsG5
0Eo9m6C0dfzVZnt0xkn1u7iS23sGAJY2r5RF0FmRGO/T8VAdO8mCWllBN1dN712V
LKSOZv7J0lvaTSjWcmxPcntytgdcQyVoYdX01rOUmjM3ZqEKdD8SOut2FLdcq/v4
7Zx1Rgo0kz+AQEi0DxwDQYLkYdLCbca7utA0WQc/6bNA92Za6eQr669Rgjx/EqxE
dLOcsMjMuiUZjzyEEP8r/99icmcQn4OjqCyYYsw9804QmhPQcWHz8Dv4uAcPecLG
FYFXW9eMEkjQSG921IU6V7n+H1taOFLLDjwPV7R0e5MwR+A1EFt9RZxJGfpvV+Js
DIaC91PNUTGp5G5cpad8JWYE4xQWESDZq85DH6guEbQj7GtrEpFqr8NPC7ltlwea
txeI8EBrt/+YLdHtTXhyufnXUowy7bYeSHlWjwzuAyFk2BSGGOZSRbayBTggWgGV
+lRYCl6Lpa9S8rcFaEA7Im1kY+KLb6mi6YUsyaOy3WazKdxaklE8p35POIiABBo5
5nWJH9bWmDogvYSJDYx+2Q==
`protect END_PROTECTED