// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
MQ0Y/f+6WLaC49tUBwUkd67+tF8iKLZ7McdTHKYtSOIRyH1Ag5bqsGfAxAUxYFZfFa6S2ruLk+3V
Ntbqdzdwn+CQ/pJO4sb0ChUeFpT5auRu4ePpEM+U0cir72YQQSuCyRfbQIxwenGjJgnWfGUK6JK3
obJdrSAG6zGr9Qif/tPKy3s/KdTbtEoNSILlti/NqC2tRQgv9FsuscDlDYMr7AB/2bO0Wdtmcy3K
RVnvybBNv15OoB8aZ4x0EH/8INJX1oQIJY6TSfHWwhwu4l6zfoPo6mTbE87NHAxGBwbX1MCCBjLi
ya9TPLfriEnjRW1G9CU1O+gbM9WI9sbH5A6ojg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8784)
Tqga8r0ZQqlI/zy/bjtt824QeF6bSOesFzsktwSAmn+sYxIBG9dVA+EREfuNB28wjUunTp88UZ+t
N58KRga+zyUCVe8UHe0xskn72bUe3PP0uUqsRmmQI+HBEXQ2h6qqiSIuG5b9LjdVDd1mcoptHNNa
YG9TQ7KOHhLT8Jw7kxxcloNDD465SX/ilT6HjyWB+/SRP9aenVOI2Jru6RnZbvxC7bFUpQ+dG55Y
0ZRr5t0v8p8GVG535NMu9Dp1DhxxfWAxGWP6PeIGiWPq2iOz6J2IdrGgY/rv77MyV2QY62UUzeJ7
SuTjQPCQWVVy1+0ejPxb5Jp50wIMDAKxXaoQ9CriyEDrlQ5xX/UHKRM6xGe0/FZFqPcG0GrHQSIh
hlHYN0njCu3XF/U2v8l5kXQUmCQmRSu3CQzYUR4fjKhXEuuYQ+R+0O8pvCN/SPWadDMaC3WUIJeu
/6gT/2jcUpg3Ov5LiqALuxACkUL/Tg0zYFI67ejiI2Ug7LMO4OjWpm7NJ0WdM0ORVv1Ci8TGkbWw
Eo6XEIPKiuzieHzFiEOUo6WQCoWrk+nV/UH5D5f5IXOqzVfUoYtVkvOFgybnTCJKDDMap6lOHftt
/EGSk0nqQSIEeCMiuz/NZ/E9njYXUklxjpg/GgmV2VhfQWdAYzQf61wwlAYrzpphJ2B0ZXYn5/el
/R/+QyG3R5gzolDi9y41sRkm0LBDE8H1Trl4xRl52CzOBxfjSCqFPMWiUFRbqjVrV0f1tTfxMp4z
zs27I1ByQ5giNJci79gIi5dijPp7cDM3znBQb62yT2hV2hc//5WeVlbjGIGkCciD3gZSixAOl1FR
igT00vO7vujyE+39d0OIwxPf3F1T8oivn/ltTda9Bq1CR1hg1mVOQFmZ9k4qr+yP6NTBM/YjuokK
PK9wSwJusWXSfMS7dvHPHK2PMNJ8tmqpgOgLu5RvFe7+qDYji4m8Z0rh/VxnB3IKQlhESYISUt2Q
fkSiBz4yvrAWa7vxjek7cMotw02plAbHqAgh5TJYu71mO/uVgf43JuzIvkEhQmRExO0nTGfQVxwN
3slu+sFZm6ckZ80wJwYjwUZrJkH/KkEjvpCGMHA7rn9ZdpAsoTMb7c0Zur5FUKpy0VgIXMzt7IBe
qnQBS2/Z0Bb7BeIaYB2YXF/yDWR6Akyjauu+ygerMF5Bxv+aBWR/z49pCR4SGIJ7WeEGtwxIcgcL
ziFYLm26NdaToRgkuMo7tiTHsuu6LjySeF4V+mfoMK0m7wpaBtPsxG9A884YlrUxx6FYMsyXdCDa
qYaNM6lPCsMSSRGNSSyBA3NdAlYAfs8umhbFsUBImoiAdE2CR8KD4VnT63crXnpLNl6hAC3CGSZV
XG7NIz6vOND25mZQZ7QDwZA9bHaiOScnEua/q0d+2ZyNsg/+NZ4KjuwEAYVMn1hfJako2IzqnJJb
pFytnRJYW+IsYtH/bqC+zSvzi1E6DjVAD3jC2h3Usm7u4bJHRGh94T9BB3uvFSvJsIgj200aq9OV
tXPwvDhkcWjVUAKSqkpAydhiyMgLckpCzDWDdwjRZeHmxXMB2pl2wzAb7Q+8ELiRhHJs+oTnV9EE
LV5V5eKAP7HakqIT7Dou/cQc+RTpxeeJIVvxuMkKRy5e4bH9YzosOAcrGQ/RpEa1inEPj+yNr7Zd
TVFYkyz8o81ayzqjEUCLU03DBqaRfyoamQLG/bdrxbyGisGyArF64gj3BK+SscawExCGYtiPSqEp
dDMZI82wOMlN3+JtyLsUaP8IYE7haUQAjxvqDAwFjkH1MYycSjtUbsZ/u8+HrIvZx3PHAZJocFM2
Lc711Kf2aikdTT7OvmSw1Qo4wf+X32+RGSyOvGwnuaeXo+JDFiAfCXbpkBiJoLiFrHPzW0qQNfyh
Kai9O8W+tgEtpCQEyPrQQenJ3BrpU1M7xagsYz/FnF7T9+Dq3LUiyyIbox21RpGme7XOlYF+3PGV
LP3MHuZlg7xpMXxlYQQEJYf8Bhy0worZv1mugbfpj7O6kFkZAk38YDgoM+WLhF885wRMDJGq+2d9
okiMJVi9aI0dMPUdUFBl39ko9/4BWrSiHs1OTzCWsxZofT4IdsYk1aE3rPwdXvQ5OCHrs0fdJML3
ToDDMb8Un81BDXaPgBc/y/3MO4IdIaKAyA6cmRla0Vy3b2QSsjFVVkH/Gt5khdJ0QP12brBe5LX4
fT1kSzrM61iB8NQY2eTmKIhGIWgu1u+vhcm7Yv9uO4KAcuvBOdYRlU6nGX8VjE8KjES33XHOjeKo
FJiYz/jQWuLjCDIZc3jb52yVQvE8FqP2+4ejCW5u9A9aExtnGHDLCurTeX8Pj0bF+NtIa7Aq6NoW
lf+rM+R6NZwJpyKSmourC1qFrAzO2SubNWX4Sd/iR6fsAbjZzvsAg34fEMTq99rvSxiG42/Hpetc
HiWg6PpI2Wu5LBIXM9W2n71yqTdjVTO6idAToMC6XIHjFsCOwSYUJkEOcidqXKFwR+arCN7Wu8Ox
LzOYa/MFAREmRVdsZq5TTiVaHYkVjhFZwpjco9xqd7/6ZkU3TEVhC4aXIMXPIUMrmLEF7PruoJAY
Zx9Xe2R01WLunDYtPhOQ11B+CzTylK965Uwn2z76txWoFlyBQdaR6FvxzprooU8bjk4htUIMdlhS
S69Htl0psIELyGtte8KTcaL6EuH9AnVIwRYckPJZfxLFM+sG3ZVpOdWm8bMzdewIOOAcvw3h4us1
RS/zA1hM13EP4tz4fqgWviSJTKhIohZD2IMrhqPBjjWhfYZj98DRPGbM5q7FvUi5yDh4BNNyaee6
EklCcxWkO7udFkKHjOuWIjiXJ9nEFGdvQV0P5Akn5URpjP1EAZAXJwDaGpl9n0JlYigkEpUcCEvi
6LdWv/LwK9Bz9rIo6A1DHUCmIfJXK9NAJSdj6wB9arVmiIGY0Ip5KujQjVG5F9sY9TOKkmJaSngR
VqEM4GeJyYyK45/pRGfwG0GuB/HDRcCMqeFFWylNLn5nFnoKA/UtC5tP64ZvmbQ7SRvHxea5helR
r0iGQ3Xv1UELL30UhCAQ2sMC27koa2AKZ5UzEe+8i0JqNBzZlHP+KR7ZDAY3moKaRBMrzpoCwUeD
iB+1/TufqCJnX+QqxazsysQIKk5jhsPq2qUr2MGRz9mgyzkLknMoFQKeI0/sCigrclwDQco9fxHw
fxQxPbOQpbXYIcwUurfSnBgMxboNlSj/AeyBf5JXb5elKulwc2sIP1yPYXX4gO01C/EqA4btkbEt
CjA2uvbEoOdBCtuDLR6eB3+uvpSwo4kPs/ZNwwatqzKbs8b8rP6FwoMDMTglo4fxjEhAVbiR2rTj
tqKxTB6INCC0d0MDrKDXgjUmySSFPvKn7Ywf1xhTHwpYtYMfNn8K+i2gzuZM0KrFAkHo+z2pfkhz
Cx+ctazVoGnmSEp9yVfV5nD0bDClizzo2mO7/WOE9tFmYe36zUbhh+GJI5a8imEYkNiSi7CYPjWG
fXk83zkIR6o7XbER9iAlT1O0ENGthIemi5x83PO+KWe8pH5UNVZwRGx1tLYR7yYlEgIDkKFddn2J
vOEUxk+15aOs1BmYWtteVgrI/AvZVLxyMGKaQoDhGbPhYjFNztFzeDA0sVyz6UvyztCUudUGNhd3
xFJ4k92omgFF3EeCHTr4OPli8CzR4SvvFa5XpsMAF/CuFaJVO43somw2HbwYPk6Wu8bTaA5hGNtV
Hl2fEQ/u2j0nB/1YO1h1nDFneWeAqEvy0EWTk9vGV7eTXT3goWSnqNAn6oUSRVHWmybjo91DNu7V
X+vZo+CkihFJdTvRl9W2zqVSlBw/OxkXvHTPW5BlcNq/DFPx87g27FNKWaD8mwhSGcczw2aC6vt1
Q9cUmcLCQcRFqRVLtRj29LUQsdgS7Pj83neVo/0JodO0JP2mgJfNPT/QSWqzm9HO+3+ZwUggOHx3
5eKEpOrI7OjJVDO8Y/WJk5vONtAEtNYxxk1o6/DBYR/aAxkN+KfxWWGCBt1EytZl+0tbgzr2PT7p
QcBCO0qltQbIAyd30gIP7dZxllFwZxzx9WSZ2pj8d0NC+JPpjvKGkJChi63KlDtlLjZnIO33ZsH2
ZvRRp3mTGGKiK564tZnOIQmrCzCkG0TtwNl7jLOqF8SFS3LBo1MZe+GNGjmqqr3vlluFstDvdRab
vE/Wi4G/x6rY7GOqNojXkWbx6d3pU1BWYZLzy5mMCx4nNCmKNNizMDEtO5/bW/G6dwFnDNHnTpt7
fqy56kscNgXNlfA7pBI9cP6sBtULFNCbeirgQijv0i6MCABLK3B6GqyRwdl5xr85giuxtvbLRsP0
GalNpDYHEFRTvszTEY+l2xFRZ5JDNoy5SW4PsgDb3YqoJYiLwLOfovabKI/5mUJjxxR6OnnzSSXC
wkoeMHbC10cQatZlavIyhy2mkityqfr2p6YtSOOS9zATZ4MfpRBxqF7Aop4F8UBVdBlHTPvzIYtL
5fFa8RgBjVnYjPBfHV62rjED4CgF43KY8II/I+4Q7YU4kA0dZ5rdWDT/WibxlT98tsexbkReYk6v
LhdEnNDG2DC1CI+n8fOMro5T/YWLpIp51lS0y0JDLiscGO8jSfzZ1H0rIHlm4gGcag7ECVU2Udbl
UD6dS7j7KF7jCkhtVyDT3An/EY9gKYpUyYuoP8Ls+V2O7XGrz6Ti3/zWTsY3gHIjP1vmUf1jBldn
5iaX/heR4Q525n9gWLLhXGeaIhDmd+UV6UYO79fj0juhWY5XDG8OlkC0X9OTobmBnNjnxix6Sb5W
Vvq/Ngwi7UzB9r+heZzFaw0S6wz6K6gpAEph5bwUJvqeIKrRcMuR02GAOsosBTCfNILSxiaZnLgf
h9WOINAFsVObpyKNe1z2dL9aX5bDSKm40dd6wHDxKSe2uGIwzD6X0tKl7sG5Dh6g9xnEwyLKmCy0
nXMm00T+YteFMLrcknk0kBIlX1ekLVHmZmd2x4IWKLNp6sPaOsLdid6AfTWcoGpTfXWoj4bJ3Xk3
IbvMY53+n0hAFOaerd4susatgq5VPMxkHtmYx2AIZP1F5ZITWjx2YOxsQD/7Vqw4Eni+8ryws84R
15OnQt/zo56sxg7tFiaMJryeCDpOKZTnAAlH0+fdfc5uJeg6Ikk6ikG3U8AqOBvn5M1U6quPECRe
oGxeK458Mm6vGNUMCcjBhuVOptg2xzOrrwCsqGHRBxR8RSqfr6r2FYXJCcNRdJop1bmQDYgukWQH
lUWJN6D1Tk6H7ozp2ZCP33Du5J9GjVlBUhyqO0dJ99B/9dbDdW3W161hFWz5Gxpe6V8D0qnNEYzt
n7ckXs3Hd2bLLTHvSXOQy1E99GeEl4qGkLWEwaakAOkFgGK/Y0TFU4e79KvsiyOAxp002NjaSrOP
XWESL3opNH+jgvSslEZzheWrhc5MsVfujhdxhTBwL23D1AJo9UamAXQz1EJ1IsHWkJ4SmOFvigMK
7y/XA5Lvsy9pMLv5O34IBbfLLm9QviDmB1i/ydcMR5IZWh3Uioy79LmUfdl8NkMn2XKWlybxFdM5
2ye69p8MjtWx/Ul7E3s7MHdbt2GSKe/8j7w+PlmJgE2GBu5bW+mj1vDAtW96rCQeJf+DzLLR6h8o
3+NrbMSKiVi5yGsJH50CLv/VMkL2RpesZMCVam9xaNrki9E7R8YVc0pvzhxMs/G/RyMgv+QuFVL6
Ml+3sMbQbdgFlKB7wX0mgihMuw6klILGoJMbhB1NfLdP9Ij6YFAEE/b734lSPMUlZwxYL9Htkam0
c/X1VfEP43mUxB0P7REWNGh3FwbVWBn6P9D36eIpTh9EIewnN+knSjA8kPgAC59rHidz0DT8Gbmy
ilqaGYS0N6U3UMcd+M+VfonWMO+SIrAeWAJtel27ceJ4J7WhzV+0BSv0F2pOKn5gTYI6mXIwB33g
/DOPhMstxNU8zL47S+dZKLsyUxOOHc1wtJRpInOM7+ywfIfQYegch9sHq9lKnNMLUcaAXiyFGSRb
VvMDpK4kDvqCnZwb8jsEK5uwMOatMviTEQJv+MA2XLm978po1ICOI9a9PSPe4+cYFalk6JCJMxRQ
YqnBmw6CEIzOfzPX5OQvKpd/ZOOWUhVscqVweKXuEQSt66UQdclHiEax4eAzElgSM6jsQedoo8oz
cDB58iXt1a3NFBHcEKV1KlcJatvRT1yHY79k3mBf/SBJKqSuOf7u8bunDJLZmPYS+otwNnNn5Saq
V5i5Fcy8CIjtlLPUGJdWEvPVNfYVHWyIf6kegDjt5Eo9jFVO285Pm/CA5Dg9AdB2QxJzQd2IB69U
DRNSjRq72zJgzdbUlqkpFhCgPj6teLhwdeVbbUTX30xZ5eB43/iDKGNAAzxu/J6fc0zUzQSGXJA6
gHjsE01z25462nxyuyvhj42phLHKZJsh0GTpASrLwqeRetYltwVgJcQHqjODc+PAqUorVOUV/Hq3
aZrTHqQ2Y351+6SYAgarT89JKy/DdW23fwVESwUo1ldIgixDpowh6Lmykat+TAE2N9BtItrLDYD3
p8g7Z8pnU4l0CgVfmnYwGT2ryiX8Pz3EnVdybu2A6UGzjY110rjccnC/mP43moej4Is+oLWqlTgH
04x5KIHBtC5jW6iUeSt9D5azvofvTN49vWbLSnqAGSq91OAWx/6AIaZdgB+GDMr7yIVbfyBafVXH
10Zt3XJHVWH8P560qVbHOBr5Xvve5rI11TN9pHBfL9At/Kcav6wJlscf8ETH+RQMPnu7DXzdX2zJ
NCO2/ZB4GJ8l+hkAOEPl0CrnqHg4YxMo7UUqhxprVePdr1otYr+JWwzxg1brBEkXQKBsfN/qRCA9
b9irM8BSS5GrSrl6eaYhjC122uULl9eEbDj9+tOvyUXbDl/uAAoCQ8h5uR3r3TlhfMR3iCKnTkkL
S5Jov1f3MwU521UaISlkq9dBQTtbt42ribTsQR0larzVbECE1/R3NZW/KJI1S8dKEoT4lmmPYJfP
kYgurXLsXZXOE2NUoo9U89Fal0OELVjK9orZuhsN6HAvVS/tnOnHJRsqbkuX5huV9PqxBKMM6uR0
vWRNvNWmErga+dze6NZY3szXP/guOy6DQTUM7JB2mGKcY+Ub5JIUkI1RbkMJ1+NRXjyadIogxllM
Z+6J5jC3ynNCulVOeehIy86y8FyFQxGelwnsXmTtf1cTrp4SAYjLWbHkFRPw5ZFdNDm/SzyZg8us
MOsvblb4TH+0/SxTa0miWri58LwhJaasRURzkqcZJbHvfCbkXtKh62ZSx29AVOb9LqgpWGhTM+WA
OzlQukQq81FW5yuE60iCiirZ++w3BdccBnVI0ygYg274WOleUcHXkbguovyvEoL+MZP1PKuSU5yp
mG5JA2wiIxSHv4NteEgOpQzg9ynJUgDW3f12dRKuNAEWyP6h6yJ26YAUihbJ94CXkYk1P+tmrU2L
RDSRRh19I5uVCf5xny6BB898GCn3ITucH11uemNGkKFvH7DL7Ca8OXVuTgC8C6Bc3BEO8Xhf4MPV
pMjcnQevVOzM6ddkZEhJgsHdsRtW6/Sb2+V5nYxCjwSgN1GiTNZmilVSIaGz+wSVn8o0jTxw5Zcc
lW2uTBeUa+kcFY7GYABPE/54HEANdXr5KzFI3X2jMcx4ElAZNiV2mWUo6jdSLk0aFfefS4/EWCtH
SVkGEmSydZQd2Pam1g+vEMaRwga1XwX/wiMacrcJzeDVNnaBoMwFcV3fcbspUikDW+rVJRtDEhNv
wcHgSG48aEFbzjXDpy89tRp7GCJ4Z1iBKbTIYH9LPdOiYpCKgcutY+wNPOc5lP7jq8363estFwE8
Jm10sh6fmLFy2kR2KbP+IfTOfSW4rk6PbR33lnQAIRPMuu0xo4GZkdCpC4hz+ya2+d/GQ2E4YDCn
Z0uNap1/yw0GsktOuv49+qiVbgkodkvtno2/eq37bai28NU7az9w/i9AuK6nt1WUa//b6bad67FO
uxG70GjNPcxIDTS2kY+uiU1IuUE5+EfZ77HDAoPZncGGxOniDHIg+Cp0mfcSeKaiihpRM3meWffX
Ap08f0O66TlBXcidY1TVpcgAuruU2HgHnFvtD//IOAuQaWW/TG4ve9lk+fxYVmItwIUVA3G6yX6K
K03+ld6acgSKXiCrdNB/3TaeORKSpd5uJHXs/BB6A/2EolQXJCOIXcnf1aerXImpNVFD1+n+wG6P
kfca8QufvotOX6yJ/6aBb24KikKA4yInnfWgN5bdDw3Ua0qh/DhP+hKCAH6oixVfYn8hteeTEhDP
LcPmejpKFm3EBr+Xyfe3NwKZB4NmVGudEOUtNIdcV+RLxU9vyn39zT5u8mykMemev6+cHbsTRXF0
X9FPKQ6Ok5KjdyTr5ib+pl3b4uTbg1Y5/PKiN4Nt4C/5wS1hn5USRiw3vrITMS2hx5VP/aeyT/CA
Q4U1tP/spW50xlOW66InFz4cEmZ1MmuFD+sjajqyjgNuKtHL0DyN6+1954pP2qAoQ4HOAa86K2Eu
o5nLKKbyqdptHbTWGtMJfEbii89Y2rIdpc/QKXYeTd55vcaiGZiJyKBF0ZY5knoUEaetb4fxfDBw
E4o8C7rC+XUNEtFCLluZOFcP7NhCUIpFUyQ2Jq/UsdBdLQn/0EtOoMnjvXmhijqf1h7yGfebITWm
xq5kfStuxjR2dTp+IH4wT9e41aLA/5u8lNbADhbYgrLLRoPVywoKE215PRxzHrAvlSwi4XSBE9FZ
eQVLspZp63023x/6Ob1JL64bGs/04JP/Yj/dq6rVXI5nca5VYSA25sHSIkHRsOQa867cBQSnRPUx
qagDJlasjQgCrK8pImLndLNxeeYV3n0dTMhZsmIL1Qp7VXNKW9ayHqkrQGk/y4h2IUz0CUVWDOnr
PRz6zJlBO1lohtzUOpiJ+c0Z1wErw2y9iyB8l40kXIEwbrP3AzZIvyfVRC4ynqZPztY8cehk2LOj
ON91ZjeAyQ3LpcElVT2Q098wvNUIcia8NKxNrSj8PV5UDV7Cv5Xc7bIU7SfhBWDHTKMj13y5wAdq
DeV3PsMuvzBBjiGUChxOUBK4Tlsn4PlaPAYoqVwFmdT8QUde2+SMmuIERBmbnwH1nriwa/SWvfvI
LMSmJX03CyyUloyktgSxbxc/x10SnlyEH7cgq6ZOIC0Z1xzoURZ5kaAwyGwrK3RNxHpiRtgdbor9
0Bb874rDyHnajdBJaJQRcgBRiLYZr7jKF7V8erP0ZgSNKIfpR2HxMBSI4+Cl3js9qi05TtpIYCVp
cQO3xVUjDHgswOhuHMVSZQeB4sVpeOc1VEDwCXr9mRfxtNx7x5u3LNDq+GkYaM4xLadC2kdiM2Yg
6n/c91n1SzNQ+stSHux0e/K4FFrIf+QIdDTsNdaYr6N4Pp4HnhEqCXE231Xb8HmdxDpvYOYMM+7y
vWZ8TYMTx1IleHpysPWW8aYv1zaERwfIYrzdOXXv5C/ZMm/jPuMtjeGRtfo6Yp4arBp1gHuQ2tXh
Srl/eYv1+8l5/b579LJEESlP7JOF9uEHKBowEE4qwgEA7/RdY9Z0o2nJ0crLZ7sZKPuEfOwwGg7z
XGxdTn3RBKzOUPDwRMTc7o4HFEbJ+jsmWpcsnQZo6hYFBA0jofjXih74/xQy6UE2iYt89MWBq0Yz
zuKPTEfTWjYPVUCMAZHO0+DBap6aJpf21/rhMP/+ItgLWEplR4mlMB9jw8ynSRJFKI25ub98N5ws
osgaDbCuJOezMPyc0oojfzAutwjkoDWx8VCU78IbJ/FyUo+eHtbI4olp3FJ3MlHchldlqlp3Fz15
gjgi1EukuviGVPHG6cUdRsVKAp4gzeSubPg04WiJfQTRrSV9WkJAK5cQVIEHt/Uf30rFdT4bgBX4
3FZBa2pNHaUEtQU/U50Ls0oglRLF+aY59ShhyKD4MF9nfrP/qicJYIXA9NbqHNp3gSAm1EBg4Qau
RaJk4/Ru7/bLbqJSNFRyjJKO6KnsaRsZhCCrWBUatYFEVPrrlYLRFRyf0jTpXVXcL5aFe1UtoS9I
xO53LgWWUABpeph8CGZOMZZ75a0lU0pxq0+fmBmxqt24MN4kgS/zE3MfM7xXZvLqWFaIGUj73m6q
Mo5PThdqk7Bt0+PkRLKDdR2wtM8AwQbotx2BM5dwasyfJFQs4atqTJHXNghkb3yO3tV2FteO9Kku
dGUtl5ZZt9bkg+JNyJldeiKqY3ZVYdoLBzWWmEdVTEDoeZXDbpb+nRaQLxTy2sjUgAfwLnj3PJc0
Nil1WSzLMDLJ1XdzifvEd154uqHw5/Mlzm5WXWm7OBRiiiZ4xDRxuPHZxmwXK8pgCc9BjACx+FsU
gg+Xd9brK6cSAfuW/Vum1/rIOP0IXtT0bBrhS/605XFO7ZdSsxe/xcdTobTCnLo3dOqC8A8Nyzw8
WefnMLLnk2XNrUk3rqFLv/fegrdhr48DwB5EIBuLVVKbutoJLs6zst269Lq6HaFt/e7+2x1eSz8I
UppT07rrk1QiXWiqEqmL+B1t56YR5LT+Xv2z1H9khNqge+MD9fJ69xPIppRtM9B4/X+MoGRhEorx
yCKBAc+qtbYET51MUN0wh+r6EmqrD/gxqV9gYPB8p5nnRyYM8mI0Oc15cDEe4L64kE+0cWjPuBuY
eJNcz8Ij8B3i+bh1m0cfTNgwJQq+OklDcUe50+G74HC3h1D9VvtAq0Ekp8k5sQsLMn7KD4k+MM0j
JZVXsmH5Vp0ae24fWA+R6qsTCnRRtNYKB+3Xh/q9z1CXgNEajKsKMKL7s5PfZ8tJgwYk++mfMylH
oUsLJhCR9x4NaPFL2d+TEcLYFXE2y9auxYO0Ct8fy/Q/wEacHt3P1Or/cGayiWtYxNQVVY4L1WLL
K8vcf7b+l1myeOikQYnUCS7XKT3sjKP5EWv9/6FWhHo2FcgKLv/wxthbUKjLsawfUUpYFOrIBwk7
faLB2PWQf6ToxUl9KLKrvSahKZJR1LoG6JU9loF7Q2yojR7RJ51L3DBfTMQeHrn6QXwXlO4Z0QBJ
ZjzWQ/rG85h1UiiU67uJmhCiOQ6wVnz0QsUaeVNMzdUkjKy78douDWFhxm52qsyHxpFt4LxRsNrW
MECGHRNY5LkG6Z9SsxW+7PJvibYE8hgG6Uyhro6Q0d8hvHvRnHteluD++UwimVtY24ty4hKxSZ8G
DGaNbMqFMNpqcLOtcjr0SedTE0n6nARerangnXZqnN9VVDTFpQSY8YfnKQt84WfpeSsGEqX9+txn
htwB+sL9sN06C3lu9ZdPxC67AgSI6/mNZ1gwfJ482n6NSFpFuB8eZaiL5SpCUmqgQsBmdIk/b/nT
GOdb4KPdbxCCsljncLCepcyo7pnnetWFT1WCp0O3JxN3jVcpaIq+JFgVqy5NX4yz5W2TW61fpkLa
fB/hI+vWe8him1tBw7Ro67boSMWLH6yM7zV/LctWFJzran86nwQ28FMiGb3ZcgdpNOQZ+/Ntk+id
T1m5AgCn85g/TU0AiDraGi5H0S4tnC9AdO5Uc/VLFsgY6qk/El9K2ZcQ6jYyOXo7UU+Jmy+Vh/po
zbP39Fcx0SsWHQ9TmpaIWAY1vJYuhiw6noK4EVxxgWtuGcrJfiP36Db9VBJfwRj//WKSpzkwiDyy
NYgGBj8gsmzyM/hRIhIS4XHIEsbqS+MfPxBrUcE8St/tbf8rgZ3m4uJEAfP5PuaJe3CyurZ4++Ku
3N+XlkSE
`pragma protect end_protected
