-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
XoFTRrI8M8lIPga4Tesgf6AtYvb87mspmwLmJzL0koM4oZTNLAHhAGP0Uwv+tPVMzH2cersLTZA/
mFM5tEtDxik91fM31vxGiqjkdfNrtDiuTqUBIGRwW0vrLPXeZQA0UpbrkEZR/0jEv5L3kAEguFHc
CdQ1ciTH8oELLyrcan4TkYArTYmE4g9pQuLLYQrjGxYTb9D1BveMqOICF4VtvRjsoWVlc09RbjrO
6x/a90uicizZfmR9VOFlMpoO0fGKO2y1BqjeNoAgM8lmS0OBSuExvuIwBf8xCyS8a8uBAaZzfLQc
AYDLslNTb5qzFDxXr7YhXjEkpa9+76K9TZcdjw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7104)
`protect data_block
NBk/+Oh5d+5KjhkhShS0Wqyqx57BR+aOV1yyoH+tD8YxUTwrYlGTtinEYaXLrRoKANQq3Qm1nW9c
M6/TS+n73drQN9W9mRGnepzyJZENM7t6QqU9nfarckdMXon5gYGRAL+AKIci1WE+HbSy5b5dwYOu
p7930il2V4jUXM+XV0Qt/myZl7q2Wke0KGphPIciFgt6O8mSJdUs5Je4oMfOnqBbaC2iLibk2RlD
JuhfO4DJ+UWhDQTUZx1C7GFzXaUbB9TvzCyiX+BSMO/YJ7ko+Wc5CzaJuolYJN983IBmEyugr662
mK+P2iRxpZjQOKltggbr1YJOIfUrLYibJNafs+92+HAd54TBeZ+2wzJtSKLzl/UGi/bMGQ3wdBFK
SgWI5G2Vvp9X8xgXjzm7XmViwuqbjTSNFEuzCfW7MQypq8iBjgV59sPvd4+c4niFG+0wWj7xWsOl
GJG5VTvHE/42oFX0aoilLGIF4K44GlStPeXcl4Op1tdgNJU426NFwDtUtf8SXbvRuIDGy/NeU0gP
49h7bZlcwtYB1N3gcWeq6VfPVDozJTpTubkWiaBb0/o5iENdZU2MaPWDAI45s+uDui5vNQxCpCc0
mTr2e7jJfBpCNnmTosMJZCCXaPddfO3yWCM+le/7ZwL2nKOsPQW6t5hHaU9AV/PD5xcnimLnnFHF
VQx7xNAA7KiJ5MrWzWu2JTt38ZjjRXbfKMSrQ54tZki6Jo8oOp+5gY/E/mNLRpIZimAn585M0suZ
3PTWK8pXNhvV/KbMzDNka7/UHMiS9m9ePBuXQPvgI+RsA05KrQxrnr1r6jHrfZtPD+sZO9wTXwD4
alsvjWp7Tkm0VtBs+ifoYghzt1wYt4xvpt2YbewvFZ16D+eHCNkoxcLeCfjiACsHeePvgMZgA2QP
1eccXt9z+RnCm2dh+lZJ6VX1fbuNwlrcKNplgUnwBXQPINCMHbaxS4FVCo27HWL9+5HWnQtZHKLz
QqmKefJxbo67Wz9BJo0BYN8re+hsUgeF8O/nSEMWr99nxsMKCtr/M/wSEJ40L21/sQoH+FeGUoIZ
AMEIUKV4/MhyH2M9L/APNBMUs71tpqrsyZd7a9V3WpHeaM+QZjVLg8lYg71sx1KLgAD85vsWc7yL
GVZK1Lrx4d3E6a9sYjbPJaX63+zLJxTRaKf8wOJ0BqThgaO9orRubvQL0tJeiCbmS7NCCC/Wt8Mv
Kvwn79u/bKVFbHhShzdhVpm5WKu60XiNiAJOqCyKEpkWRZXicr/0DU47ZxTPENs/b+dz3rGwu765
0opfF/jqmFPSuLSsCLuJovLaD/E9GBWOMFtzrw5F1VuzBRb796xGm4CgYC7ODUncrqUsIOR3OZrd
J/mCQT9ohZQloS2JlyxUZIrI/RuP4e/o54dNcJXXOMUkeQLyS9gf4Hf8+hjWMMCRO8t+550u1IlV
nLqmrFKpTdQIrNVmA/61GvZvoN9bwdoojENrcZgehYvXkUSSe+W1yWaRI63IbFPgIPRmwE4ZtmSY
mCLr9HmZqyAwr9UpRe5wGrXQzR3YoC/ftss+u7lHrOgMI3lTOzzRpnqATYacVnR6AgqgLiZ7QioC
zYw25qaD7lONLjMc1tybYNYhDDsZ3Y2X0tA9N0waWeUY2XU6h0/eCPwfDuTLR2UJvHHrVcZl2GZ7
Ga/1L6WyssDpWl7DMMoxdw8O6zt/WOX8CHENCiLGZcVXbDJ+EkRKg+CVFo29lBloc108g9/dGNg9
yostjCZHGMF6BTjHINKClgkLWz74eTXV6TzHs8Ie31CzPLs2jqaquk7+oakJWXGiW0MdgEnU17hj
/oXIV/5QtH1JaNwBZ3PaVDPSRPnGsoHSLKhbf4knG4mO1gnrGWX3DYLDpPqN4FDyd8lsttfxfS6x
a1Cc5GBq2a2u5tDsbvm+9YBl2aNTNQmQC/Pn/VwHkbBL3N/VTKL0biKW5XVLUZ067RAniSK7U2CQ
bt83tHtK9RTD/UwrSlopVjsd6TnCeG5ZtOpxAA3veLOk5y8vioOEpcv9s/7Yisy1yoH08XHIktAm
pAiKmC9XmjX2bkvUG4Io4lkNueJiy85kjyiWnnWcGRLaUQ9Vw2WnM927OyL7Yptbyblkds5tOry6
KKFliwQTvOLMeBDVnmmdSKWzTvJ+P/VkhWRxqNpbUsEPdAWoL2YDTpfGj+MD2Y6EfJvJZmHjYlda
WmF7MjiV7ZtYZN0EGXgz/mRhAnVcfiuppSOOfGo8sFWkM+q4mSDWkx5mIeIx87vrEBzCmXebFHiD
pEx2WVBoi/8TMcf4KrnnpUjl0CB1XP+32L+4VqC75hPgBGuSy21UzYhL2jqhrBbPwqRTFKY6KjeX
ZSd+2EgYmAB3kwuGo/I+YESE+XyGV4MrCPy64oS2HwXw08Hni5wXY2w08YtpR+BRqZRBMu1pSuqB
4zjv8Pu5FOhJSx7UqMLOQJfXCiM5GEgG/s7z7f1NZH2t3BNorntYEzlaMKPienwkUztPYKIClaDo
QMxZ4i3/ej8EViGg0XgIkwy+w1ISv0sdk9nNjTAPOSySAuZ/EOtqJ3TzGwcS1zqiaIhhI/iAkI1k
tChItZSzoroYMeahLtcyL6DzvrOVaPmsQ6moB4bfrq7tXIPgOfdft5GIdMEkADz2bbRBPwiWVnwJ
cAwrPUzxkHRK57/1OUEXbBhySv1Dhw+IlAF7QvwAwesanG3YwW6WXZhCzN+g5Mi24EjGe0nb500+
/dp7+lBG1M+XI4jurOnxqBxeLZDleHxkiVvO7XLP3TV0z8ca1GV02f5AGKpFOQqBlGySj+VlOFLY
Y9Bu007+A/kKl23N5H+vW+3HbN+MwORndTE9D/vKDZu0bLEMiQo7WDQxygZfFh2wzzLZuDccYTZi
4ibnGGo7VSc958cCjU7aUb0sYeX2i838wHab2ctz7Tl4q/dWUQeBzQeabLIfBeLNM7l/lKZ8bA9F
v5DECLSCF5XFAx/nhh4jK6OKN9Ds4cK6IB/lCX3CPAaUJp9y10JR7NmufmqznP/126156qpECIjE
7dUJ1RbhgV6/fU7hRqlYZKEnVjE8tRkijPSm0m5COhKmhCo69Uk1y2+UfqBpbTz/tFI2H/JDwWp4
LIj7WiOMIOjz3vSEmIuEGYiTUeLsMHgA/P9n5Nv3tOyNKtord1/wYAeolj9feuV2s+94a5Q9A4lM
pkenzI2UYSO6UhdCKJ4MZQPL4LSti8fDUw34XRU2/WoxnuqQTzzv30yldk0anZogpGV6MYUpBAbu
7SEYh7E5sKCGFyKAjO1r7EJobJcqlwZox2uU/WPgHFESfPgX2GxJLd0VmieQspYKf6i4S+q95l3d
PFo11Bsei6aWQmHzGISGPmHSn4ZVZvjY+5Fsa479kxF7LVvzi/5gqvDsn6UG+omhzB4pViDpEBkg
OZ4QIg+PBV8/d3KQhu3vRa5Q/a9Vuty2lDlDi3xpW/qKJfmQ11ae/KJ0CwZm/oL5PTwjka4hNWKX
nXe8ALH4yqbPHWgyfW/2iZq7Elb6/+6WyqHYCiDpUDm2J+qzrQRP6lShdJ4hyblV1G9Yo5adv3Wf
ZvAeF8J2yZjaC5xouCSNxI4Y8/d96e86CSfXlYu2KkzzcsO02OjV/smlTkeKbxn3/6DqCdg8Djsl
4S0YP9PDIM8aB4Yve+Tqtd3t8ioswhie7gwCEAzSWhhP1A7h9MLhM6AAUC/XBshUnYpuFpdFSFRO
jActOhuL2gP2Fufxe3A9zz6G/UDOmBKt7eBvaqgIyrsy4Z8NBKPCNdHNEQSiaefsubBL7fMn1sLk
yyujoKx/eLcAe/9XTWeVfLTDslI7AcExIXTVyWO71BL7Hlh+qM29EhVDV3zrRJxSHWTVt2TAez6/
32MpLQcJjxu41lHyT7YasXZunLeyJk/VgI5HK/pUfCw+hpt2G1lZRa/oeprI2Sgq/Gu8OgihGyHr
6Fw4cl9mV3TYwkAyrTKlnh6DqHDip29YPGFh9cHjNafGDbQVJCL782ZUsyCyiztjTmtX0NxFjUFS
EkZlfs988Cks2WbZ/xI+HjvM9FWCPWLZDrw4l0kmYE0kKEgqEkJrmHj34Rm70QZgu+7DthziOFjk
iwp+6nxF/Q9AZl1Auj52F9k5HQO2JvE9b2fh2+YPjpT7PbWXCFRVjeRFMQb0auvezmKACVx2TXTa
755Od05J2YGqL09jKnbfUrGb52E+IfKrY8ZRlU8ujcWmp0NcH18mPzMRsx39OLSYnPuquTSZPfYZ
VmaugfL1K5Md8cV/1aIAtJymlyCIvWzmCxVFRzABlSNASnxeu7RQzYdJmV7zghrwzcupLC0Vq5JZ
J9M9l020GidI6n61mxhjfw2nIjrPdyGRaSYQl4n8ayXe6q3SP21sKUzFoPyCWfxuC/612n9irx+J
T14+EeOFWE+Hdx7luWogcw9UJke9SYd2iu/PgNLJoqyj7PnvLpmlc594MHzYzpxvags2qJSHWR2u
zm0a48zVXPul9RL/foRM7b3+UbOhMGDYiOSk6sjhlSaitq0yXpBoi+1a0swH2mA2wWJp8NwnsD2l
wwljEdE0+rZ2aT5SecbOpTDbAlRKUg13VOj7VogPnS8/aM8UhlclEEkAJiavDTDtyHwHinvV+mZA
mI4LEkIDekP2WS0OD3AMWYdQK/NEZcBRzgtGsBJiG2QyjR6OBC9VjvQ1Vr5m7U9RKldxaqw1Vfa5
DB+5VQpyZPqzHPexyARHtUeMPemmyk60rzYoUnFkkbbr3BP34aYbbW/VJOA10E7tlYqkc6ZfFTeR
AUXseC/Y3kXxqWbmzQ5zS7NwMgNyGNIX/ZiruE00ZIncORGK59enKvt4zl2jzurCYNZ0cA23N7Az
1/R1LWD2FX63sOon8xSG0/VQzyQ3CSpXKpx9xtuoz8pjtzR0jckGhCi/yFkqd1TXgJS/o55qmiTg
25vdgTKhEjksI1zZDz1e4qp+xjTJvt41KkJoFQ+txgNLC/kBVnfR/w21HJsy7/NIf7VK4LzJ3OXe
zvHbk+o4xfmGG0WZgNjb3VhpEuXwsfvhOuJ4rmvoebrNSDaMUq69nhg+mECo6RWD1R6qnwQGztzm
MOXEYJKbV9uHqgSL/xe15SPTwXftNz0c4fQFYUN27Vp41n0lkXklRXd8GYFUWw0gUIiXjv/rnsPm
6cSMkQ/GGCWCGAoih1g48uHA84gf5P3BVBAYH2FGeluFfrnZZ6aimFJwY2/WMWNbjW5FAN6qzLDC
qU/Iub0rWwhVQTOtMTtNs3n4Ha0EAVNMHW/iD1HmSHl3kLIUAgMILos4NjMviZq1vejtJivZb6Iz
KZx9f7yj+OB/5xehG/t0y8xThZ1FpIHysvAb6OuCuVCkWbbORafwsDJg9hhXXGyvQKZHt2TmrF3l
FFlBnFe3XYNsPxw86HnDDnfN64pglhBiMu8qpxL3jrw0D4keC99J2ABzn663RssB310TNGboX+5v
uTox8YRF1N4cqqqLuINlOiiIaABciGGm47a8FqemCHJeKnPajrRiRdjH7Gxfts3m/cUEOz8I7ip0
ymyrzp7xB/YzDwkUpoFY+5TRd6G/iEscUCAHCMxh2lnFjKPqu80fkeiogWWazMM1125xfXPhBlSS
ME5s8RfcbEgIuMTsYLEei1iGTV6Ijn7sDWGr04pQvqTx7P4jkw6nd+HbDiv2Fbnk++jQ14qgKioX
KEDAaUGxsygpLzHpxziV2yKjebTtbMd+hYzcWZwYoTJvtH0BmqXWpf8/Dc64C/rlErWGTxp8UZNK
TcuNhCekPl+V8QyI4CqiuXIf82e8T+wwAxhNUnbW7auOrKSsIDQd8dpySYhM7cTzVWuffbW4MuTP
qiHSOK/hI3dfvEeXOZ51YnmYUtUfHW9HhncGUOZL0ZbthBpC5qnXxr7YX6uex1tZfqz/AqTOj8w2
n1yec98WZcim0bzp0pQ7tEm+d7Vsx67RByClKBmoVyPBte4yay1Z8nUjiD40FuHiau0aHhrCIBlC
w8R9SDpPDdPQx0ksDulnAobFGTkDMLVAx9heUoVuTU02EeT4KqL8Ub+JIkXsFQSUjLoqBdyZn0ei
G0m7NnDEftdfu6DE+kvSVk99YxpkrZWV9FFfzYefNUsCNR5EU7ejdjBfFFkW+tsTAXg/Yt79b2aQ
sd1k3SNz+YTdaYJZTxlSXSBsZAx53Pc6T5txMqdfMm4Kr2Gh3clyBBiYJaZUMXXJWXqy1eFcaOWT
fSH9SpWrVkLJF/7iFPs0AuG+HjVOTyefiIKvcx/R/jqS2hjmDUGQ/FEdUkgbWziZ/gknqT2ucQDH
JCmhVLC8GjsvlW498VGrfzRRiUzPdjxvxKMInPNKVRZqUFH3KSkJhSDCH+/rKqpgGbGHrr32h4Mt
Pllv4JX2/iaesEqCflo8tz43m+9I3JxP8P+tSqPBX7nKTO188SsY81gKJvFKZRHJTLu+c+M+HtEv
xQJJry0K4aamIlEK7rYhjQt4uvs16QRQE3AYpGRk2FWz2QsT0hxaFH0JGKilAKwY19Lb0sq80iDp
2x6ogS92ZbIXjm8C11Ce9nrPWqWQOg15c5Dg3L1vTnb2CwUXYLt8Le7HEXMs3LLuVavXP4C2g5vL
mlFEqJmnD8U0Y2hubBGVLJk5Ob3F0FVW2qXoZOB8xB875Eardq3j205vYpoJUnlLQewAsZI0Sk3A
fHiNGOG814cX3Shegonk/Z+2gMCL0UEmqGzBzGkS4oD3Hd3nuI7mgRBFyqlp9eoCpEY3s5J9hMrR
/ZL+hcK7KDFYWKEQFRk4hHfg2+WwvUSIryB/ABBoA9/m2OjrHagUB5oBrstBJ1zjkCYXs4Eim0q4
F4CPgPk+tPztgPC+pe8wttOV5itk5nCbUzExpdpSK6Uwcd9FQST27smE7lPte7ZyVxSiqDjx8G19
hl9Fl6UZ55uPJNpc/2ab/Rat9DEB6V3HUcutvjMgBrPz537srhIRrmTbs//tEWHnYJ6Bw1ACvbIg
VS3sxC0xh3BaJvbW7VYJM5EdLjky5jbY4op1d0WX5LdRtTBBu3Oh51bkeCvBxl2bAsUqi2kCCUwr
eJAdkHmBJ6s6bHgiaD5233yShu6qKxvEyb48tLvuP7otAY5U/2WuN9TkpJ6WmXns2NQcY84lB7kw
cAY6eCEQXTpFn7cZB9qeSYq2z8chz9JqPYdJshN9EtoCgTrxsJuEzhAJAZa1LgJhbzzNj5ugKKJe
WORp8AQso4nb+gRbv3TZP5SC7EzDmlrt0kwtHFw84BbaaSImU8h4u+LYUh0SOIWP4Z9S7hU6wdgq
WEnWShFo5yV8B+xhQMTxDGZ6diOssVkyIFo2hQCIRxei5wyzAGagGGXODViSM96HSfqpUJQCYmev
X8DV6BEaFL/k4cl302qeA8dEC0jqmPO8csKpSmmeBSWBclZjrOX7kg0z+Yi6GOnuG58yA7DEA0x4
jal+QzPgobhhYFLqP6wsIZ4plSdowitCVnHW+M0BmLc/Ji7e3/YPHuInyYWU1L48N3lWLCP/zYQs
RpPnPi4nvJnIvWqxdG3bYY5u++quWcNiuWZBa3xzbahInOMjZxBet8f91QWGe3hGlJtNr5lYKJJ8
ADxkx/wT3XCTApMHszEX2m9QKvs9F0iUjupLLuI4nsffL39+xaecB1SI0yjHdwfs+rxNgRiGXZfg
cm9F0aORjdhTrzbWpgmN9CwmfyMZkXy/mfN2jhwoXujfoCbbiGZ2HEGTcXSWcj1PfSkmp6bRvZwk
agLM+uK1IDiMb13FOmZWogREFqs0F72oaA64BWhXkJr2ALUl3ktCa4O0vdHSVrJ9LXOHZ0GGFam5
a6yzUAcQjT3+T9lT9yqVN4FctoGZ3VKsQOv9ubV+HUbWj28cYV3ZEkRn+hgsA8a6e0+HoS4am4Gf
YDyGVgBIzcJfvtaZfg4hc7PFVrdiygc6/HU0i4OTCmltlyFUiZReftJz8s1qyFEUSMtjaTloHWjP
j9nqQWItoPWYkIdhRazlzSv8SnrqxyMP3+I5U70QBEnsow4pn7UkaXTRipF3WSW7Rzk+GhmHVKEr
iBaAY87c9ra4eyc19bZZTGQFGpSrKgim/YnwBVAWh4eEd+iqvr9eG0kj6WyexMiRi4JJz/DgOa5k
JW296Ul3lVxVHphUt9ijr6NjZBypZsl3N/+f1CGcWNU/PV6plaUtf5+hNgeWKw8sSsWbQ5o1wkAF
EJGPC1bs24K6bFt4PYcfQ3rTvg/jMsrAEJSVG3NEJfCRJrSeN1kG7w1+LgD8wMNYaNsJQnlA6LGE
c3GjpEZ4VGMRCgoMG1jWn9JRymo1GK7wj3h9q5TDjZj+abAlWt5MKDln5T4LxJYMjpW1yIem/r+I
HcokjvDqrvQfxKJSqSEjT7tYhKpQlBZy564qHrl9zOsHMKiB2DUd01kqDvD548Cmqpenw3X6DPaV
guhYESGTuTqM5d9/DlcMk4PgUbw6NdkkytUElJKOB02VDsbOQnJkm1HUZjWiBWyVczPJ76p9G+ai
NZOeY0jaqZQc74fvhunXG7sYlV+nu9/Im2h5oUNBwn69rtWyRjUUV+FBkFEfXIu2JQswE0CUk4P/
Wq65Iot8HovBTIhjSwp+8Ozmm/7zHYIujd/fZI0ZjSOJ2GE6UOa2G4dWJHnXSNoPQ740k2Si3Tqv
XJaOjpM/vhwB1RiStNF2YF1G8KM3enWF0tqN8B+OfY+MXLvksGIFZDr7LbWLcdtoJW5MyW1lz61D
2fo2MIVGmQoYECYT7vZMVfd+RdHwfuS0t1aaxLWiu/mjdSAOQqRaDX64AFjF6igR8zBrlXfKnoKY
md3p6VGgwe+e/svdoMg/eEvBBzEo7oTPXEJayho2q1jcuuUcUW1h+LnolxHcIGcpm/A521A2WCXd
PG34voWTRuEbnzCQc4eQXhn9ONqtZLaRg8gE28Ofk3d6pIaSvi+V6l8AWqbRE5f9wuufTewlptgZ
eKNP2g1ioy0M2GuD7dXtMsZO5omXTp2y4jKjLeX9I1Y4XCPDaG8M3XhmrqdoFVvmnks6VGKUb0E8
2q2q61R21j1aWTHXiWMbqfnsB59Jz83h4ubvRNyhMyQhtCyPbTfn+GAYIn7mDUIYe7yc+ShZXs9Z
WeRw2IBWhld+jfXGLVPitV/km8LuvmIR+PjepUaigeoOXHQRwa2iKNN0qzvYhx/dPH0Y+6BmyBVK
koYUWoKK+0CH9Y3Nmmko4YWNzpcFwEe9ZxYdAW2iouBqXRi7ttNy/IDvZYSu4Y+yD1llwZESNAVy
XLNQhDdj50Z2iYjp9ZujrOoRWO/q7G2gVlCjltxtrBzjWOPq6fHQ05SgtnMAjCOrDKnFlkkQkklm
WX3yQohMo0zy7bp4uE2VNrr+VQxb5kQ7tHJh12R9c/Amk5m5gFdjpikoTz7DhvCVZK867lR98bOq
rDIKxYYDClVU8uYgmw9fqyn70OPBV0kZbSDHk81QVJpqYK95
`protect end_protected
