// beamforming_delay_calc.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module beamforming_delay_calc (
		input  wire       areset, // areset.reset
		input  wire       clk,    //    clk.clk
		output wire [1:0] q,      //      q.q
		output wire [2:0] r,      //      r.r
		input  wire [7:0] x,      //      x.x
		input  wire [7:0] y       //      y.y
	);

	beamforming_delay_calc_CORDIC_0 cordic_0 (
		.clk    (clk),    //    clk.clk
		.areset (areset), // areset.reset
		.x      (x),      //      x.x
		.y      (y),      //      y.y
		.q      (q),      //      q.q
		.r      (r)       //      r.r
	);

endmodule
