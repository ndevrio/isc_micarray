// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
HQx0rBlgrams4YEH6/5A6pzRXxHH3/ttZikUVTuxzvjQczTjASr/SqGN/9QtYzBw
jjAebf4dgqddJzH4HU9b3Dedvu88jrMgai8MfaDTMKwpA4/D6C7BkEUMawNGjEzu
CpdmK95nFVly0neDjy/dvTDhrCW3sBgaR8rj0jpve4zLj8WlTn1GBw==
//pragma protect end_key_block
//pragma protect digest_block
sWxSow1HuRzk7fXpLb5cbIBoAQU=
//pragma protect end_digest_block
//pragma protect data_block
F3TEnctKz6sLLh1/3sby925x2kE/Ja9RHSNxUsMlz82IjgC5dYZ3DrC6w0O6iHR2
Qkrj6aSjiRdR4n8exZavYyXvPKCSNIM3XtXujYXgSPX4dFYsgc40jRG+k6boI1kw
VuTbdkjSnR6TWi0z38L4Pr9tZcY0b72oXDR5zRrnyczzfp86bd1uMQrvZEKjofS6
g5lW1Xq9r3ZXpkj6UT+7lk11xKxjBNhiBPzoBnvSldH6Nfv7urF1ZRPzTRNxKQua
KQ1ecEiuGmPw0NndSeK/IdoZ5DKHxkJSX+2jFkyleWCiytug8a1MLW6iQm4kTFRb
aGoTUNeqe+ZzD4o0PXodYXeTA8ErgqVfTHr7bOC1N931NNa0S+bvZCIfVXNS2Ejo
xAemTGQ3quv2wbAuefqT+0IY+Qub6lhVoB+r/WBMHj0p6pplEQ/NjNCFxtyi1CCi
mYsD2EMb6ydRWpnsIIgVgNBr/awOumSfCaBTLkIL6EsY9pYahhYNXhrJ7N4HLVEO
6ACbAALzTG+1Qyuq3eMRDxcbPFn5cHYLDKLcgp8wh6D3KFPhej61QNZfNbh/uhvd
CAMGOTigSF9BoG4lRo+Sn7EcLkayCvC48Cipu8VnqtWEcCERFh7brhS3SoGUSiNc
mN7Usysk2CfbGk+J+DiI5TGa80ux8Ow/e+Zka8BgODIKFnZfDanM3cN2Rw8l+Aqb
1GjBhrR0eKR/tavctp0gtkzAvEqkmj81OXkuBCgraRheB2MaCIHY+XP00DPOtt1K
S/qtleUNXD1jVTQgzYXwOEMT57oiW67BNZTGv2WrcluDJL4MZVA7XwvRWa8SCTqQ
xL+qb5TXJ5OwOm9kmyGRUHzpj1oWGxlON4t/zSQQmlXXzBq494iSd8ev3C4QN09a
6L8NQcZ6DCKUUy+nXcEvPmjmJ8mCk1+yQ+00Ai7CwiiKoxdZuOGOB5jufzDTYn+O
QnLHGdl+DP/ELXrqJubdXktbSE+UAEJcnlw5pXUCk6A5DTpj8A6TwDW81bMnUD2P
2LrKmYslnkLMZ0an3SwdlTFU47mNQvnhXUeJz6rwBmNd8Chmt0fLiOiJuDdB4v/g
s8tO6sKJrQ95vNiUITx6BaDHyTGDnGpDzowm7aOuWlwpYgMgmifYaO4qRIcBoAY7
sylhU80uQzQ5dg/rf9LG2J2ZwUYhu9RbMlvwuAJ8xc794PQmITPK5boK+w40KVuR
MBqjy5y182p6ily0JqaNrY4BKKAvVkuna5nQDVf7zmFZrLRep5hc21dLfDyYSFBh
h0J+NRdIbv8+Vv1y/e9RKjjn3VfPucjceysopHHIkOdQuz/3DAj2Mnj8Nd+G+8yF
SjcFmv2HEEZHzezjjR1U9py5p/gN2aVOQIbBKLCntM+3Eeu6H1O3t7J6sTQwAmVc
xhqaPjh7xylxbSKn7y3PYHUQx8dN10F8Z3UqAKokr2hT0GzXpC8QR9oH/DmIeJdX
Za6e0L9ZwiIeDyYjU7xWfyPj0hHAXhRfUGwzBwLx8UJxFnz0jk5dUDZQACsd7UCG
qVbpu4MdbQYVjQU2xt/UlqseZvMNhK4ytLq0iKgTQ4REkCW6rwrwgCkpo5gFpqAS
09NqKvUd4GZRWha9MZhLXdJxGH7o6qbNZmkyXs+NyvapXFj5Xu2XOArlj4Ap8hO7
l7H6n4uTvadoCSDafwCdGPthD1rawnfyMFKL0ZPOpJzJmmCXCwKi74umETzpZxv7
7chIa8xxj9n1Lm1gpE3RavqKMErG+hKjTi9xKbEqTtNtO8vz5LMXvoeUyertP0ud
zn77Ns4BNEyjMlZXej6cpnsK8Ddpf6RNPZcu8hwC//2bPzbOe4Pa5Lya7X6HzsuX
WkG9sW+hguntHJWflNYypufb1YMJxfz8J0ZzIm1kRaUvKcjdoz+nKaRdKxGwZA7M
d2hcQUirp8SqdLjywPic8rdT/+Evv038Oc0eWDMHmOnIoIH/JWMKqzdIkq+ua3Ae
UkH6E17b7tJV0ezUSY4TWKJ9SioD/3HijziZpAB0S0Kh9AdbLQqmz0DY3VHqiXF3
AN2hCPaLhMWfkTUznal2XiFGHm/XQ2kBnpkvFqx2erPt+36F1ftqalHOjTpUZ5ei
FqfR2ULdis7RXnJfpjiSopF7JxRfYpI3lHGkrjIaQ9FFqIf/NiOFYyuImI0SU+e7
G71/ND3d5XwllQF7ekaMRfNhl1WnnD7RnpoEuLDDhws5INpMxRx2i5VXyr1tWgYa
XBnIWLJSwIIvolJIFzmk1vhNiSJ/U1vQALtHznoBa0a6kHcTH6QCVpTELIYb4YdG
KWknQj5L8MW77OVFgag6zkhDYXDWV1qwuoETVyh1Qg/YN89zi3WkvHOMlwV7VuFk
tNjcoZ40jU2/Up3IsGWFER62TeRh5kVEfZR7Z7MvpGJ+BZb/SKZVFP2l/dj/Gss0
W223jdZSzFjV9U4grslY4b6zzWt6M9ilgZMtbCpltItGufNF+FG2kiwfbhWI4PRE
HdHQ44VNOHkZvjcznBkeYjzvXgkD+CKMRUF8yLMfv6ARUrGX86xdaKUBgultMjDt
jCIi+J8XszweD2eeC7JEfew7aeG25HThDNS802KbJ+KGa1SHK9plxo7WHBfsHfiP
Eh5qM5Yvv+K2VnN8/wxf1QcwOzkIxotwYhCcLjokIJKT9KKO+EqYX12NTmCyq2z1
59g32KsCnfg7yvQ9YYRlt5TN+1EaEkyYc7YnEFzOAMCDKWCydZ9OejDXWEAqGQrR
YOjl1zS3y7q9Ah/9+qjUnA7dbs4OUQ7M6okLxSupDDZxIHEbeE4RKQqvhDIAnfwz
4V752BzLYgc27xQgVd6Y0bBJxkF6y4SVBkBGThEaku4uui+xrmnxHD3FUK6qRsaJ
62BXNJFh4erfR/wjoP8UdgPb/R9eyB6a8VVdyob8yOhw4m0gOQT9C3Cn4qXXltrs
XPoTYrAIW1KywJal3wYgqO43IsXrZluYsEN2MR41OV9GnEx+nLTT5Y3Nx1NDBO7O
TK9Yf5YhTvZe1n9ra2hiHZGqOFMVFvN1gMFOXxZD5BUc49Efu/mzZTZW80Y+Uo/g
aZaAwtgyeM+wzjceXRJOkl5NoD2nfAXJ2XC8TphLbzDgvlblyOZbtC1Q3Q+R4Oxm
PVkEVbdRn64WAMJCxy+ULnzF3wO8zsyFFOh82IUm52eH2zPVBgmqTfI29uIrB0ed
DN6RScC5PI+W2EZbuATQ2AM4RDj5pWBMztvuRx3gAheZuCPhmPA+WbZxP9x1l4jK
FR4gGbSwehTsoPiL4uid9vm6RAdYiDtmdL89qKZlwJgfkbwcFeGe4AN4k/6+/Ak4
QPfoke3J//DoZ4nvJHG70igxROSFvraPv7NwJnDV9QJcyv09wGz1lcLMJvCkZDAj
ill7ufTWPld9caThPNz8qpOtmX+SOwiEOgkyNNGEueDyBXhnJxQZXayFrpo5IBfi
pLNsbk8DDSup6iH3ACUkcC8F6udEu7T19/j4youtDqRvBP9aeUJeVgthEkuayVUi
5vlRHYLjLgX72pdlYk9EDrBJhFexYlBeVxEj2UKhKuDSBq7nq7KgfyadUHPsQY9K
fMj41myMGe8Hd2K8lrc4U2JtJlq/GQFWMtfZC6JdwEkJKCyftP730mavq7NblKGx
0kX6sB1RdagPH/5rUxqqLyK+kDSlacfhfAQn2YmwVQH1sqvTbTjXwqRsw3RHWaoP
IrxKmJHan3JRsRMQtM1IHLWXM/Y/h8vVaJ2Cjp6IRsHezCtjRCxfitWh1f5fdFjz
2nLhl6yZt2Fgkb+e/SCQ+7EH+YjNkyHe5XT1r5tBmdwooLyAW1FUrl9uuXs382I8
Ug30PbQbmdrXkYpHRkA07bO4ekW/oMuJEcS9CQpt0ALu1uhqXHpNb4xxDp9u/axF
V6RkV4FKMH2gN/hMs8FerEzGXW2pc5nSeZ8E0TJdj0a+lSyLgtgcIOFkzKaviwxI
2YDolFeMZf1kvSuY/D87EZATSPefxw9aH1qvRvf7fR0JC2QIIkFRsAwXQDG2Oeu2
uPhnLYMEYn0+RUUZgdrrDEbcmdKIEdubQoHCXb88wOjIIc+/A0T045aApy75ycDl
Cm0YveFds3JOI3b5Si/bai9sWeGn11HwzZKrDhPleVhwPtrzBJTDfRGv7zzV3fkv
6fGkPA3dtOfvaX6MYbaL0gOqcDV6jTUXsgu+qRgjU1FL5wWcSfcHKAzmidp6zj/f
IskWidQUeENulYh4QbS+MYAVnTqB7nr3CDmcSG1BPF3AJmWrTYmTi2ISU8LUCFOt
dLflYXonf2scj3zxpJwVNnqno+NryCgYvYhTi2L+Zkg7QFqOOVsW3VoJAMNp2wUS
UJ4ih0/7c2sORvdvW6SgX1cCaHjZnrWuvGs9A8mlUue3W3Fy/S93VOheXMOYI9LH
e9uqpeKwVvPazIRyXRj7LktjmV0OnJ1Nkx70szJ9wYd5f5aTTZ7UclfptpIDW/G3
fO9mA4S2f3gEAVIniAfrhTproFKKysmWimWAYj46ku08uc/iEC4OrGjWXQcoK3qg
ng3iLRk/958zjJjKacYSewRKmvrEeUWUtBmT/ElSsRlfXpNc2pJm0Iol5pH7VtlW
72Wqd9sL0qz/JNHDSfrbyJRaQGGIdY/hsMbRsrfj9Q5Lr2v43n9Fbi5cOdrv8gCu
ngF6xpPjHZTedn4RT+yplHY3UXeKY1SlJsek0BUnfiHNxytAIkj9omSFKaJusQje
xmZxSHBhabGksxsSOgUFJWlfnmKneEUwfz6IQEYljDLser3NRY2hxNXcC4w86IA+
VnGoXk3Er4IqXiNZdRKQcvQyTTHnbX06zZmyziJSCHtQdBoS9y8EL7FMSo77CWev
Vvl6pVftbmnlxeEt+9wjocKtTnQGLR40W7Vh14r1BdzHrmMeHgq6TPChVXUMzleB
5Cc5T4/VriXEp7ju+4VnmuIp53QZrQLPR0szqZHAi6i/5+5w5BbMPo1439MBf46x
g8OoNuD3NAj+Viv+49q+mRYCnqHYoX9eGP9NKBdAoX1mLPpoxwKExi1sCcAOAnHu
xW8UYZkaKS72Gc1XKyBcAoLG9NpBlXsg88XsVjYuFtb8gduJe2JWUCsm0ofSvzt9
nwMFGeHF2h/imN0HRsldtAFfBNmjzwKdEDsSh6Jzd2BJddG+CBRwIuVSbSPS0I/K
hsUEUBOHph8VL5B7NVZ6ChmxNep0CfcTUXCPN5AysqWsrYMa+sIxCVqff1lORdsA
IpyCOqiMkd2AnoQSNPvVx4GUgMO036vwEgt2CiFG7CzUnbqR4F7kWxL/zcjxI+Pq
Huo7QyHerTljk6KJ70DaEVlVfU5syA85HfKldG+fAi85YDtiTEH5IZBw23paGQ9I
3elXnBf7yjzuo4WQIXMQSqMkl8aunVVr4+esr1Gok21Jon102r7fRPHX9b9DYb1B
2JWXxLynImQswHKpyX9N+AMZgwEuBD2zDne8h/ZCzVBojbsWBDTYSDl+b95YLT7d
x0dmjESyfHMkkIHIcOd0duNhYS0p9DFAZrC1B0gz/Ra2c9sM9ScmDctsyTIf34e6
3BnjhpV236HTWSuNALH3N+EprZwOddocC0elh1jSlJ7e0PxvobPN930Q1+ybK4Kg
Z8G8qiiy6qJhKakv0UTZIhctqQW2WgWcm3x/LNyx8TupCbznw3x3O3MdqK3Gu+zS
rzCnlkAaUfri6NqEu3CgM9uIll5d3LinnXC6qwhwpdSREUgQbnOnKUbhJ+MZ1zmZ
HHPjRIytiwfNd4agP5cZvb1x7pNcc8pLur7ixazunXmslym/wBS3KJnjec9nOSAj
oV8qh9AqXGfZOwfv5btWnNHWn0GYz7wrkI27kHrYTPpLfKwmffVgcwKGLmnQLVa9
NJcpBdaR9FkYt6PA8aNFdPHVOY4WpB+Td1UG6SrUVUeBGXv8qzD7Cq1MXCsowLHx
dEs7DaMR+y0RJT8JC9RvzKtrxCq1jgNYIAUSv4deg9X2vihGOo8M+9I+hkHfEqZP
s8XiLvITZgXSavEoU/0eetgVPOPId6WMLdR6zGEC4f0pyOxiiBDVFayRVLo3GsC/
I2JSh2t9KV99mHDtE86j0HW6foepxdQOqBc35NXqufs7tmvtC8JsP/cAQ0nLGkIY
lWtQfQxTmNT+6jJDbz6lQ8JzyHnR+VePghQlLHuJ5AK6Rf0zv+2XeEkqAxFYuGSF
8hxE8dD8abUsd0iYvX4slF8Jyj2Pbl72bI/Ervb4uRATeUchDq/de0vXUUdh7EbG
T0nypxcI8MgDqSNvLMtZ3nJ/KbJe6CrdaCL7tD7HT+PwVngH0Gsqi3CNI5lkHAmI
b74J6KLJPBamGASl4PGlqJTMD1GksGGjEH56B0Ls7B3lmJ1aBX2avByZXWM6Gsin
LE+eFymSM9/10AoJl95bKyBscobkTdtjeZGMHYoP+OjIxQuTznGkBL5Tc1Z0WTi7
KoAC8ni2h9pDTPMZQ0swb7YruGdi5Hp7akWgaRd+I8BcnLZ5Ggb1xtmisVD+Hl0e
0yQAONTtIUedDMWI0BExtg8I3hBMTg+fmE0quM/eplxqRhnO9/vACL7ASUJeI9iD
eLba672SO2cBwFyRYFoAmUpMp8Ax/vXApqfhaoRAb974pscQKjpEmTAFQf9XOETS
wfCM/8A5VXONEpdSgtuCRZ4HEBjlxRGYyUn3PQKnaWu83MVxg+BEcEkdU/b0Ek6r
ocSr3TXvz13nlVtbnJIJZrvYtGMRBdjM2GIaXVePRgtKSpJmAi0/hhqSivd9Z/xJ
kwlPTi8/uvTzr/iV+WlpxsAok66zf8ZLWSLPFPw4Cv3lbkJPfsrt9Yg3F8MipQDL
/pBVeQT56+nVpC6BATztMkrRfbzFUs/KuS4/GR0L2lMG6IJM/Bv4pJXvCqpTH1ja
bXChwBokLwgbOIKl56VY5b6s447w0zGX+cQCp6yakzbRXrqbLBVHNHHAIx31LwC/
0yTCP0ffuXhX+yBw0jwDokBOj8w89U0bGGRQBnRNqfcRdej10fWNpE1LU8afQY/H
hIoQokWD1eU6J3E120jYb41QIndeSpcDt68RBDxxgpisVHJd8KiqOEd9dFnYhuqX
GigjpUTYfpd6UI7pmwO7J7CaEl2Kb2PDTch6zbcRa332PLYz1hR2eIN8qw+SCJD5
0M79/actuLHGFk1zCKYBOZ4299ISJedKK/Gf+T8+uhkQLTAAv8KM7nJOW+dRsGKO
F6EQRjfhAPLmV66jlpKkqxrlD1yDs2xQYIRWxRdbWIChvPuC6NtQh+i89Ni7QZPv
z2bbDtOUG8MJb/Yik60DBZwlxoomJGRXWQDf/jBkaLk3UtjIwtANIn9DDS3MQn5f
GmyCt8rJN7kbDWAqLUGVI6oryv6hKmL5T2/eKy/Afka0uG+jow1VYF4VDQ7lrqq/
Ejs4bVU69MDaRF/uCgtcWyKt1O3DTqFsPFMyYG0FUk2L9eUNPJclOmPCxKKzv9ga
apRq0KUCo9M1jX2jJrt9m/LOVoYD38NqdwzUbytJc/QSx1z8syz0N52Jg+WwWpDo
XTJk9sKGjLpEOwa3kQjq6OzI+EHad9MhKY2UPukaADYrerPABk71e9qDxXeO7JwZ
YfBk8kGRo1zqWh4JT8Q3i53OOcJwm8qBGMz+d4pdqASr585BqgT/vQmlEW/9nSO7
oEiy6nqKxFhK3gi7+VFTymOJ5j+r5zPWpFv+JDWfA5JBaz2Wkm4i74fiZknJLMbx
D/cik0IiVOfQiUzlP3HAbygf+8M/L/VJR5Ckvs2RQFMG619292l5pohxEhSEV4/o
Y2/SVK5u7bs6xXa5R5PPD2f1Ho0Q40/EKth5lcnTsYGJUMwKGisJjr/6yzFpQ7mt
pVzXm+GLjHfil/704YxWxe40jgkSMT548gg760mc9pZiChZHDXPYdeQ3v7b85t5T
EpZ9tOHUkuZb/KHoQ8ml+mWP2DfWxK27TnhXzOf9GnnWjLMUzTY3O58PoQ4OdJhd
u5zWdGiI4JD2z7A7eMvEWW86632QTNcbxB/2JB+WlfaZh/N8RgG8iKaCollUwhQx
5h17vUf9AxVo79zW85PFFv+jW94Xm2xcTcCKGYHjPg6fz9r//Xdr08jGQrqwgZO5
RX5h3M49bfMxsnUWaaYcQyUUxCQmob7cQe6ZY2xWQUxodh3hLNSpq4BA9/B/ZvdU
OPibo0PratlOLOcQ6uob57BLj3jYE1qPeA7lSShC30fyATky98VP3OVuJ5RORiiK
mw//KNtI6MO0M9UYAvDfzpfOlBmwp50zyPgdmhUVix0PeOetoZHyvsBZiFDErdux
r+EZYcWmlU1XVg0povzyKJvtWIdpYnKhq8db9aM5naONS+Apuj7UFtwuCejJXkUV
731nabEocWBa+aCBPLV85AJRjGwxDHIFjKIAsFT5owtGx87j8pozFjNQzMc1jgvq
l5s65xn6ZI+KTOADTGeDr4SOauFmLAKud+a1Fo95EXFb53Rxj+F/XsZa1z3WXALk
D1Llkwc4Ps9x133IhfjU2MVzZPzeNOwtXvhdSFT2E1Byp+VSDEeczbSHGbit71ag
gYeyyLNmVfZMX4WKg6akDa4zBLhU91k7vcS6pth7EtyQDoF30PeCnICfjYE+05F5
W2IXf/ayN73Lcw3n4OJfvspO2W3lo9ko3ZAUo0LGxsZ1j+/ma1iNEQLgtQcO9lgz
LJg/5ucMOqgTRVuIu5hX+C/YMvW5jb8lFSGUP+J3EP3dmyEHIvSZw/t4xmkpblq4
2gA0xLdWtBWM/4b3ZKKJue03CFgYV8agFk+QDZvk96J54ulopoCnu3u8zPzB94Lh
IoC+0q2cXErB5NbhPDna2eJ4WB4yAhCcQpbL/QrdjQHtQDuHfTNhB0Px/VBlCsyv
YdB3chpCL34dhHU55DiCfthopvO+LN20reIRNnGwV+1TiYAMtTMIY4mft0L++99Y
GUHOlwS9s1xi0+EAyC5qwLFI8RVLAolmcs6PV8fMoOo+rMjrHr7GJPuK179uuqG7
zyJDfjinr7nswbfGb1eoUsVCiuN74yGs+XGF46Tmfe1zfz1ENZBkSRZaUoKsK/ac
HRkDLgVG96NBV6jNBdxTCtUCxrtJk+Tnts+zsLOYiVHHJTp+mSAO3OFSzSG85NAI
aqj/D3Kb5L9hhSVfg97nWRfmKT7tYgRKBWYKr7KDvqZmFQFBSt9vNFaYyfR/Eu+h
uAzPeM+490SvWNmPr3KFtkSOFY1+PSz3WWKuh2Bj5ZOlEVDPS/v+YB8Bh69pAK44
W1+TKN36Hc4WgaBIZ++MWP7YYih5H7Tl9gvh+/LzrmiJvjPCblJWZ2NT7xMp/AV+
eBqsWOnarwTXTNprD4VBdN+UKdnMXKXxmgmvpZTodhw1IgBkA0tmBv3yxBlS2Siv
RtScnjy6ltPoFF7fGq6X+1y+VHw69W8cPGegmtdxhe5bh6HuEOQppINyy1gv7BXc
q59vR6CAROnnR2AJnFf7GD4dmY576hclmYEvQfxdJiGG+QEKu/x41TOLr+SquYnp
6s4B83HBcNCtavXWgU0TxybSRqk0zk2NWxaASQ+mK8PmEOhQaxy0ifadlv5KoTRI
4vFy5Xy//h5Ln+FSoiF+xtSY3bzX0/u7ji3jlsy3oztgwrf3VKe+HXJ4wdQ0lZEW
qZQOQnLnR1SYRarcj5hGd39HZZDCgpA6ihhzx/NFYqw2C4QJvTDvZvkbTKg/NoaK
VPgrD2mVOdVDQrhXkFwDGScJYmGf0VnNap4z4h9O9PM7PtSqZcLvw/5y6SA89ub7
Pwm69ZGHzmXx3tM83TRO8O70NQFmarVgQ9z1GKP3wSDdhAzZcbGnLMQU/YNiMTeg
1Nd089EmvDSVXeJAJfTAaOaHdet2UEv64qYXyUB8uus7ExxDaronMYnNQHVPW7Hu
Os2V4NZxsOqNQ5HR3ERWFngvh3cP83/F3dBEhxSyIweYwxUfY0xLvVIf+6tvxnwg
WkFrXsqevOTyzTv8GAstETAdE54U6Y8X+ZGwOSbcfYJfCOE4Q7h1Js9bHbpR1bwh
mFnchhy16xI0y3zaLUvexm49LwGYuOK6QocU4PnGH+aJ6K65L/RuCyl/SCO++iTO
l84sOnjSFyTzTSUbloNLUox0hAZoQNjDdD6JTv4MLfGdDyghzfQLZEb7y5P+/HDd
onki+5JBo7AF2GON/5+pKk8KpDk/h4trQmfuBIM/X73Eul25IGErTFAIXL01BlOq
WcNzAN9JQWuD/4qIwwxK46Q91ezdqDm2Cd0sHoR33eMYjBB1mO3BbcMTgAfvMNPA
B6M8xR4nBadSyqSSbSlQb7Rno5OO6YNGwk87FAOwiz0/72HiztntUP0NJhN2mipG
UERFM+1bqilPXfrZNm23qB7Sp9pNTFSNO1ozbl9Z6/MSkgI+ZV3Rvf4P7nR9k5Ry
ZrjP5iPFbbPp8en+dnrkRFlaG3ONeC8hGr5X7mvgeh6SDph+UUycAtVdZodVAHzp
mk+YlrGeNH/wuY3tiozEELHefdCgkl5uM8Jz8hxXILmdpxMggHPzHlhM/N5I352h
RAr/qmzI6X51XzEXnbKdr0WycUqfh8ju33iWMKY0Q7osOn2l7iIQBVmutXu17T99
c24u/Ju5EUjz3cWZ4UeUIGDHWJSpMjbig+p/NTieOSauQdcE0YIqWLnK/v/5LA53
uromHSIWNsVIkN7A9sRGL9XgFv/G1QLIzr+rnrY4qQgwH7UrgxLu73VqfwS/SiRq
MC4ah6pXqfDpD22/hUUqpd+s1WY68gwUA6eLLYpzLcQD3AV+LnhV6pg693Vv7uBi
Y4HspQD4etjvZDmSv52nCtsf2bRBEJit4lIt+8G0V/isDXxOpjpVw6MkZO6/LncF
7H0pWUjS+/V9nCuPvSeNvukocqVrkkVX3zZxWkPfggAJxel/pq0qqQsA6zOtGOD5
6rHm7d4dbmROih6rsgLSeM8LkBAZipwLsOv0gvNljMRymBjYQiH9YXvX2jPLBpzc
EsfVZfTeFL4DZhbAnD2kTkeW3pCH3boD5oTEXAXMbx0lXhS/IR0ot8LDErQz5pKV
UmYTo7gE5grK+SFbXgldCe+iU4Wc0ehC9lfhojnEkG1H2xxSa9rAI3xFzxvFfRi0
WC4B65wvFIPAoXV0puagQLHGj3CWYDSmy7GIVh0KiAcXKQ0ZjMSNUzY2fFifssta
BL+xpdutPlw62Ro4okkw1NtMlY3IJ0SGQZw0RTW6qhnRRRu/JvpSmAEYfBvZMlYW
v0WaHUo8fMcfIkOKmCuYJ/3tbu3bEMgb1eQMfP8SEmd5uijNCUswDabSy+T2PTDL
lryJqkmgRWgZCzmnq/9orGBwj08OE0YE55uYd5o+R+fsyaQrGH81nfPjqdF491yL
WmbrpxGbR4BJZdn0mNvKmHwEBLpeoqxd5SbY0yDQ8fac9R+xewtN/3RwQdAytcf0
zQPEyAOo3F2kgWYozj5P6X8ko2+p0bCfUwhP45LgaGFhb/g9AZZov6GPxfE0V7h/
ejAh57EunLphs57rtF20AbcQxuOo9+fPQSBMuZSY35EszRSx0SHdKqBrwlGNzsDY
EPPu9jX5jo+fLhZlwwYGCwIzLv32L5lmgl96Zw43ipCFMhK7bQsfVsrlmXJelDWJ
5wRreyDUmWJ4rTCZyxHhcA+hVMy/KOYWU6W0s/ZopYrC5DyxMBdQFEdNqc/Py9mv
Zmpsvv4LZ2IkpndZ0KC39SVNJWx0ptxdS8+r6xNpX2PxEdLUEmzNiPFB/8+fxkF7
0pr+6cAbCS5lYW9DSgkSzCKgJxopTOnPbeoSpR7DpAlzQ5Julfsly2p7SNnAPIvl
JuPtq47AKZC4XTSd7LcC0vgBrmod4NQUCYwP+jxH3Yo/kO9wmdY//aB9vWF699C/
3wELrm5dZYBlLE0DFhbCoroS8MtT9658Cxa35geQUVXdqTEUBRdNDwyaSO1TrjWs
WaUhJ+OxJYjlV8PlA4LlYNEUt5lbYdSIgd7h22Futx1jxYyIcM7uOkPuA0qJu1Xw
BuLQ4naArRrD/+v9A+pfuq3hg9Hvrgwm3Gyb/QgY13YHVZOHgBXU9AQc1j50okkp
EsCIGIF1bEd/A3ZVWcTRstcGCWGI/ZD2ON3uICD7ZkgLFQl3fDVlKuueN+kAhPs/
rLoGbyktY/4bgYNECZVr5RWdg1NMtPTGLG9G9pJKELleVuugvyDdBhiYWMsOt2Fz
qNOKTha22pqHr+cqrAZvE68CnfwG/OmnfVeG30+dW7CA+UtjKrCPX+Xy7oyS/1eX
CBcrqUFX5VOs19KgrJrXtrBrTxj5OOJ+u0kJPF0hqut26lxgki5dhVesjQGL1Mj0
KeLVqTIqoJxxkgXTmHVXVvvni3B9zNr3LRvab+D7RuHqlmhVyRe8V55EGfyG/55O
n16HG355SlAZEVdz1PrCt3pBQtvF0Zm8xL7ur9bIUWrlYN4LiAaIXAbshNTsUF9L
YE4/u1Xrr/A284jTC8/f19MPZYh7jrrbJiEy7jnpWfjgBZiZm9BCtfIdxhHFQ1xR
qC395M1HE6S7b3LKMRQIf9W+TC4Epfiwf+UVdDJyWKsGN68t11QB63xPMaMENc8r
2xAhjCWM0/23mTlbLFmkJ4Z3FmGD8SRA3UACP6UGprtmiwKI/THlNkqs0oteaqtt
FJEy3kE3Cqtgz2T5f5UnOA9z0BhNR71W7XCBil8lT+4g8ICOgCLMbQESw6Dujymm
U14Q7Qy5doZ5CpnBGeR1FCPTD303ab5iLVbjjKrRPercx2ygfpQf2ed62s0FUlrQ
tYhO69DSkIJcJm5RFw/WthzSfMriZ47f8EvaPLxHFajUj/1QhdKRH/+kNTBcMcN+
eCXYg9EgoLcqlJ+q2UkJuo2dBc0ZTVRdSfRxWIujpoE0CdHcPK7uywaNucL8Y8eg
y8RTDTRH49tyiyiC9Dfq5DO8NPLk+sIRdVRK/SLkH1HFbjXdaqkLlLCgGzjnO2qP
Q78xt6lWNGZZEUytlfnbwlEEBpoKesfgVYn+eKV5zSCjLLkeyNeQreebh22K0ulf
qLBsC+srjn6Ikltr5v/4u4cvjmrSZpa8B8SIqlLi3obJUszM9GJ3zvfgrK9pXarM
Xm4uzkB8iJuSEw7CEHvqXmY8Ne43gmJ4XXzgskmeGMp1Jw4FiBdeWDQOwkicE7C4
EvMhqrhO82IevgVephD1QuZ3TWqvh8c4QDpbQFSp9c9IT4w7n0VlBIFbHtbJ93xy
2p0eRW4twXYNlkRyhwXzMsT8Xj82bTZmSqK46DPDrHBG2D6TQDHaYdt+1+2+2kWK
BwocI2lba8irFoztrtuM9BIwfHBmrqJPTw4oXLXaAXaYeOy/hLe2t03KE1ylgQ7L
vJDKZaYgYY73p4cGA7ay2ItoeeXjtCB20+1imRK6GsGeeAxBMhIkqb/uQJhs6vxy
g4N2HxxhavZooObWklOF56ansHo6mmD9RxQXJy1KarXKFYVDUVYPN86wMU0T3ThG
kCObyOl8AxoIuvqvqZokbaWMW0x6qj99vH7ZIrLquKJz9qrajdC0a6nlsAt90woK
oGU3Rw6Yps6803bhmeOSKCxrl9bm/DscQHNni3Tm9/zWM3cXuvGsijBmXpmr44IX
OFidKQdiE9FQFB/br4gmF5KhyqvSjCiKM2hQsm+yMXGV5gr26HVhdw2k9XJmZoKv
47eeJKIABfV2025mZOb8yJydhXxVLx7ZERsacYNqL2RJQnq67RNd6RZk/uKwJyg0
NNmuA5mrl8HrXJBNSqzYI9GWJmm+uocdAD5nq4Xxn+TYgRgIJiOEgCTyXNpecBRr
UgbxCAQ/gJJkBusIowPIxPGRUHrPobnjosFMtdsu9gsXvaXdvkKWFjFZdAmvu9Ty
GqBMpkfAyTUXt5i74J2B3SyaXpKYcYzf+CmIJzqRsYPBvkM+AWU6lBALYkhr8VcI
UXma04LxTh27p1JXe+DTitIdT2RO412CkBjnWkwZlRN/2hWmYFaxfVbPi024izMQ
D3wuptaHhEgdILSYnx+xythuQxFuaOUP735bcS8NzSi0MJph7yCSD4jCl4Bks1xQ
4quw4OJNpjfSUBEN2tS8MR3xJ/Rzm/O0RibmPZ4ZQbbK3kKyv7/xBlRgZbMZk9wD
qmjc92hVI6ckKMihNxZlFUgXT0+OE19VriAzQSrhU7etjWkbEHzHHsqfeuKrVXx1
6G+BEIom2ySOFW5dUdZS2oWy3QQxSPouHfPB1ifD7i8q2ovsgNYO9gNkZ7+pMSQ5
cFXaJFTXOVRq66pC9ZDgB+Jq57k8flraI//XVLhzQwknqlT2r7pu9d6Z5520RyFf
YyDEYoNaW7857uvJa/VLboSWFfwP6hZ4Rfspk5uxYXgCvhyJHKDqAty7ur2pgD5S
jd3RA7lOT2yfbnLLbZLQFWIaVdm6ozmEh559AoqJ40FTT01Eby7sKXC92Hp88+Cq
lMkGcEo06cCstqxy1gpo0dr8KMB59qBDXOcM/EAq++HmdLwZjNaOmEH5NZBVJ4jn
/8t3s4gxX2kkjsYl40oC69OgkoPlHjKoHLpMaGWZ1aCs1fwa5F4i7n4noUZmzhNn
fyiNFW7a1SCXJflafCfTPuVRPS7DfDjW39LhQx64wkhKR8mx11KlKOk+P8V5rzbX
8Yk81L2R9LJL35nTwV3D8PSIbX6UbYaisb+Lr/y++YhvOai5D12XQlD+6PyQK+QV
nzdQTlq4F6lLeu8oaqtJOlLDcMUMob5Js17UBCqCq20gz0qX4yjQAxaz2CAJL54w
DwSTCZ9xEMXDjwy8jDusTiVl1RPZAev9xumMfDVaw7mn7qSq+j9frc8vdU0skmcP
ucoPTLX2BmL5pUJnmg41WfAYtSAjs8X9EG578W6tZS0XX/4aaabILAGFdj9WNtuE
/UyL1L5JBiuJdYk579ENJCVDFu1c8kFTDetXzIxeEQvXGtdwZ/F9ve3EKSNaLZo5
gubHEEoLpE1qs4yv0ZK7MwQwt1/EWxwRJ/LCX07fMhirsEfzM5KketiPzcEyFE3a
PRitvrAVS9l3nS3Z4o02DJTgPSQPFYJC8U/UOTQpZwMOKbk1md+w0svGzC3pLE4o
H4HJiuz0N5rW+asnHGGo+75nwROa+o1+sDQAW5WPWtkuP0dxTq9LWg0sqE92nwup
YW2zqTHEULV5M4OTYKWV1RaDgbkriZmHxenpsfayyb5rUBnBJB0AxnO1IRausz3a
MbzcawM+WQo6yeLqffzW/sS8pGBBOVs2NgMNDcQo8lU5QcTPZDMucCYt7YWPPyNH
wMWRbMXBiKEj1zAHP0QM61FLlwuIjIHWnyuwOj2kSTt64WBUDE6jIp7GPEB2PPlX
yGCRdShxXTRsCyiU3htNAq1LIdd7/O2oXlKDYt+PutY+q5b059DtX8gfPbFjDPQj
H1VaJwGH9KyO/iV7JFNHvJKJKi/D0Yxo3Rc+oOAnVpOip+bju4UHesxhQvUtKkpS
A/bBvBKVBpausAC7owEeXQ4A5nlE3sOSfNe45qGynfPua1YLNJITMOT5G6qwjLUo
pOpzm5R3mAdnFPsaAGUylwHa4zeuUjC43ZBetNusu1JPc2OFmYCJ04v+YbbXVzQh
ikC7Lw8C/WC4Zg/bEXMYxq+j8p5tLnck/QsZw78XoYbNwSRuDMxl4ASdZS8KFU59
LQOuvjAytRbg2SCDgE0nKXBPPp2IDMsMW+9RmJZejmOHgnp+9W5Tc8ZjRpXBDkOP
F5HIvBxKo7eMk0RmYigOKcNl9kFuULf93quf1kf8blMT128OH8xWFaap12uJ7TzU
CJjUYo0K170CvYBjbn1ZZSjOi1g9YGY7KJtb3UA088mqtWGzmQPKADA0fY/3WLGo
dkMXFtgsKnK8SZIQzzzpA0ED+X+Y0vbSl9NcfZOi6JfrcZDZXidVHNSWXnnBTZTt
pK0LOtiLXlYG3tyB79AFuEPXWMJyjMQTi4MB0wxtV6h9wEpF1dU/bQI5zBv1JhxE
n9w4qtWuuvit/OzvWd9GSA3wKK4BdxTnVhxf3pXj3mBOGOLdrOeRRWlnjeB5NpFG
B2CLtzqmPbhuEZMmQu0iSxaFdWz4rglNvppLU/ZalVX37Fs1CAxczQDlLA5ZS4Ih
hmLxLrA3p7DYR3/DkEwDnZ87tpeiDvvfSDX7NpoXjgqXpV2SYnXYbTTy54qV8JZg
b1m6GLMLl5PD6ypUhcyl3EiSvt5/VEcrbZ94NTCPbZDqph6+/RABxSgEzwmPZajJ
TxrVox0qhgW+uqhiJzuX5aCGQSVspcXIeRFdaaYGIjT6zsgJV0XEsVnypAxh3QQE
PTYxIgPmkH8W0Cnd94Dw4evX159ERXAEW3HF6Jln4+Dbq/z3QAEfg1r4NxXVGL9M
DUWs8p7ryCOUQU7hoDM/JHfO8CWfAlJgoeykEwbzDSnF0ZwJdxzabei/ZdbDduti
D2KGThOmHqjNyrF/4WLXIHpfnKLV6s34RrS+H1/7wgVWKVCyTKIgwJtIdW7/u2th
XUy07m1Gn28/2VXRBqhrjJgdsxNZnPQ7EqqmborcEPuexd9M4yKBhJXseuN2e4NX
CxRww+21vPRo692R7iIV2AySodVi8vTX1lRVYRHy42lYc+8+r5Xn1INNLaU8dl+l
GK9h/HaJwwDJKUZa78uz7a7ZgrlFtDjR4dhsVkOha679GuSh4boQ/y8LDKf6A4Bi
6APXjqzF7gUoA2W3YlWzR6qi528Q0i84LfkjivwKpv2hG5rda4uvzREcWfgMLZFf
izIm2IlUejb0osHN5u675axjvL+TUmK4tkHQrvJrr15LA23A11Fwv6ji6nkMQGJ/
b1adi0Tb+6oZW/XZEU4LwiVinONsll1DEqCht6fMWp8RHmKWokJSGdW8JBBskCGi
9ZXPo/a4eEDQdlJ3HTWpIGkrSf6LLx7lODFBcEsGYkEvRccMtOBuHU0dFFCeFwH9
9GFjt0MkQv+B7dHng2s4/8nCxJgiUawLFN48C+a1kEV7k0eCpfnkg3ZUT+1hraLd
fmFPCMNP5BHhfHPCMYdM5td8iBe0cvaTtd16twW0j3zXOJ7QqNnZXIVWqVAWm2P3
Rv3xCiLmp/Z3BWSsecs2bPHJlesd2UzewH1gzcBpN5FMnBtjHbVsBfFh9UMazZFS
g88NoAROoz1j63I0uwe+hoj8ulXXFipzDsQ/TLXHHyuLRHO8n4VACjjwpf3/l6tu
f1r/OWY0TCqaFrd2VTLQpasP5YWh/gh9bnWnLFUQ3iqUV2dq3F5QyfNqweYXE4t8
cOa1d1yx6zfhotFdiSTG4/iToJVluH3pv8TkOrZ4NATnwfiI5AAww4fEEX6FEKjn
P99FpERhbBw5sqtnY/vLZOQXWlCqIS0Lex3eq4jVhztLY6wrcdHOUI5ip8ngnlUi
+jsZqjM09oTobzeo0Qq4FeDDjGeNN4kItN/CO4vYPlSwf8Ue9tJn48ZsqjwWGuaU
Aob7w6EgEZEkLR1+Ho4BBBM7IhxoFYGSIOv75RS3YzrgdL9kyvYUacISmCtFsjQN
WhEGc+VC8jnpjmJjZ0h4cThU8Z0epjacLiAPbO9/TRb2op2FT5IQG58gq6ic3wQO
jMQwhn4eSEtGBRl8VJAy1jv7ULQXbKbTdcEb8Zoh1OADJN5v5yOY9KS5JeMS8xwr
x4cMA/IHnoOpmMMCFaPJWDZwe79Vwf+rNOQyAtXVFe+e/TgXG0QR+VXQ4+VMUCBg
e90gV1h5YNJ2Y0QWky4CnQNUrdZJtx68Ooxc8e5+/4TbZtENvw8LA865tFxsj74s
dI4sexanV/UEz1PrmKZbM0hmEW5nQC0n+sB1BHJ4udgLjTd7ZR/k7fNAf7R6R50b
JsuAuieRy1Fac760e/uNA4gK6R1GuHlI9/V9+52YAjlVQE/CScVq06MZzrnOoKdI
SDGWtAKl+3gcGTK9U/3xmZSqzJBZd/HPU9uE8g7LaPARMlyJgY83L+202RCdF9/q
2RXcQhAwXBTjwgl4hn278y5WyYhLXS4NYuuXE1PDQYngRfL0DxzkxOos9hyAYOIJ
U6ZWOWr/8Ty2KwFnkChlyaNpdW+XIQbqAk1MupMwXtKkkXCVqm/6f56kYNPac7ec
N0JJf29OKfBJcl0Ie/QBNm/S7FdFrZkrnwZfZF4dsRAFdHeKOe7qU5lI5/KemRbB
KehGDqRyadD9gZ+pcjIMOn6FVw4cZMoDzNWVmhJ+mCUH+reUm9H7TRYbGmAFM7si
0kW8HrUwPQQ/G5vU59Ch6nvbj5UKHAPU94G8Si9ePfj0NGeEe/kJfpQYBNddCB35
hrg/Sf8cKYwBbxmO1T5hohPOnTtOIAqmH0K5KG5ZT9w=
//pragma protect end_data_block
//pragma protect digest_block
zWyuX3PBQXuIyvX7mISmrfvm3Zk=
//pragma protect end_digest_block
//pragma protect end_protected
