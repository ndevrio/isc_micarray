// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
6wCakJt01BFbFRIvnwx1x1BNS+3gYYnZ0a8jyoBSGZ0FYhuplyu7E5+efIIPMD9/
FVGcyNmxaiZFwsaUW4cFkrG5xwIiJ+TAYc7D01Oau8x3FBnfaCsBcXqElfjz1u33
qBaVQwRZuMvXFR1lGEg60qPC6ydYaYtA6tz7u2Dv7F38RTAYmuF2JQ==
//pragma protect end_key_block
//pragma protect digest_block
BPbqqZ1UErTm6MAAu7RkA+Smy20=
//pragma protect end_digest_block
//pragma protect data_block
0w6fTXL8SRL6RuLG61JV5lJfABbdMuOjqGVK5lDTxH3qRsvFH9zqHDb1L5DCFZFa
t02Haib9aBba8muyDslP1sFFQaMpzZmVvd4EldxnmglnErMunmykCbP7fLlGiGv9
6OZiDmBHCgBQGj9M4W7jD5bCzuVE1IXZL/pjnjfSN7jffCU9rK5L/PaqgrM7lJbi
mhihvcbsSDsbi1us9s2U1XVEVYYHScHKjhBl00IUPQyK+48lPjhQrzAAlDSR6knz
dhdGMMBbbDmcXOcC0IP75cKziBxQ1BiQ/DIuGTRqVoJyGR4CCiJQLVjd47jKHhIi
EG7OAZtKRhSEkFMXncPzxYIiE5nzG4f3a80wu8Z8w9m4l1s5ZayTL8FZk6MUTKG8
K9lc6pLPTCqFiEPL8/zq9zzMTj45BIcbDGHhNPM7LoaBVguPe4DPYy2pS6WiLiyS
XNDQoPIaPwbuHG2yZ9XL6sCaX7PwCpW1fEj7shA5P5S4jKzfZ8peVlYemQc7iJ/H
d9lDaeF72mTQU09gJImEBusy3mELp7oCtchujbFVAZXW6aG3z71A0J+moy5QAKDY
IH296U/u52sg0xDdsnz/KHI/8BGFvuKgGXaE5NLFknQcoy4K6Ki1mmC/thBwvfmZ
EqZxcTf2oP8W7SxUUgisBJikn2vtVv+4Kx+golGEdlGYs5DdX3Ws+W6AeA+Pmiap
kXVZmpD8Y4sO1aC9kaw18t+66hIu1YYgEfbsNl4i/a7Pn0o6aqwbQpiuZ4dVI2NV
mm+ynOE5LVlB5B6tIpN4EAOBhPjDN2CPmEeVnpke/jm5XgEWcOwx+ZkKvImOowpP
5Mv8ZgVXbSk9M/fES3VNlVf7MhDNQAvNSSPRz9zMYmcWeoUdnRLme0lHp90JW6SY
4Cp/35zhhXkq2caH/4OkPBkXKkMS7aOjXCUz0AWLXtN8HI716jzt+YH0XXy92o1c
qG/+zdsiELvGkdh1TmdTe5AKLAjtsw5j5VywIsiDV/JZLOScRpHW3UuBHAIGfLsy
T6PksCJRszYu9m5xzOd7LoMBPPLzBfhRdupmoaYU1P0CSI9pahzVTpmzQN2cv/+Y
vl/11KLfchST5cbPCMC7gD2ruxOGrdwdHN/ajiEuKNni9OFfjwAmcnbwU9XqfbdA
m4XNyNUi8lpP63ES//AhPP5zooWElsuPmbsh2KSKOKnR13/3lZi4Tv1BgBRJjvPx
XObjXFncI+xgJLkX5yyg6JoPyiPX+yfp03Oh4+SkuZDoa5pnelVLBerU+1cTmhpl
E4Y71XyFiRhiA8HW98fQC91VPdpwTRxHtIrlIK1LkoHZgkfYm6q4bM2U/BlhVbwm
dC0C8oN8ovUbpfYOoB3CtcwJn+CZzdowW4jMqgIHB029mzGAWBntRso3WPHSSIRh
JN3CpJ6z++EIAPnrZVHVO0E1ls3OCN5QOQQvWyt4KRmx0V0YHFztNP9uZ6luLeM8
a8zXs36VTDkJf4oSxkfcsFsFvF2QJMkEmZmTTARnFmXesLtKz6WlwAaJR6xuY6zV
3p0ctSI2sdPiQjOS9IeN4Z22qX0teoHe2RYJograBS6RtmgbcZOfs1K7OtsfTBoP
owIMFBNIXFnJdYUAVrCJnyGwm+ue3uiO+XqFMN3YPRnlcQO9e+DvvDthz7+IH4tw
PJhoWs5mrH3fqgVQNvaIjpoxiNwQmNrpy70igudrCtD5FaBj/x5g2q4lZ7cD3YdK
8xjoMeVoeMGjyOyPBQmpwqyNRzCn9H5N2OKKz8lwxQLXH1aBcF/ZpLFdMPY4PFl2
p+mFzA35gxo2v4I1M9mQpELFAj5evXUPtqM2yg2ZmQZL3a3GXmzjQ94nOotL/4Fg
WHbt/IsKPJ6zR79juTEccCjj5ECmP3g6DZxd9nTYwlFbL8JVC01bkiuOv+rIXISt
B50dXTMTGl24/UY5e2huEqtZb7I0/I3ggZIaTiDQUCEvWXOoGsGNdLr1Mc8+eZ3y
XWDUbinp7qvFMeKeet7o2mz8TK+Srg8U/bOXn9qXG6UIdQVQEdhmSAIxsj5fMpJ5
2dWGNitXuqQ4fyeBDZQnk0XnL3GU6O+EbE2VsXNsebEt8j9wgLSZYe+roLxSDCtB
7IeotymobW79d0IBwaX27wx35xGFWRCT/6XhHsPDrWezZFg5HJ8Xp4mSA9qzK0bC
lddk/hQIk2kjF8QQRjrs+143x3y6fqEGr1H1HxgHJniCKfaNokwEJXbelVof1sVD
KU00571i+Jq05gwoh9KzmB2QAPVEiEqxj4jjFe6k+/2zBGvb3oXW21rT9o1tZDQ0
2EXFWzoUcTWVPyb6KwnRQGSoKQOjMxrlch14/1fcwHU77Jh0XIvuuCTzfWpcyc5o
miGKRBkfOI3HBP97RUmBiDDSrsqqr8YrmuegHMg5ngQJ0PkD4gBKM7kjNsDMLkgu
UeIWn/YeNKsDSuQURyUZZNsRsD2o77+oC3+eJXgl0rSNVBzBAvGwW0qqMZIJRL1+
vW5Q0ok0rm7ycqqM5Mn8JeU5L0p90gncY9Rea1yxudicBqrp5XuIVTke6OiBc/aE
UMCji3X80w2uXzsrwxkqSx0JOURWOVNn29TXXEAP79IB7RwIOPcqUf2RU2bIszw4
+60ApVwK6qHnHkSmG2yVSnK2VcvDrbigb5kNCfNt0CIXCjQDkNO8jXsiY42j+W7H
P8FP2NbCyQOexxLabulZIVb7jFQhUpymzhw1V7T498lTWW+NWHkFnUpLkB/Spumt
oEEcFzNnkIZ6HULnSdkORD4aU1Kk+d78GGauxsc98Iaxu6jnuhZ6yPh4bzWePPzr
x89qpV0iL6t2j25KFB0iKp+IYcz/Go3hwfNXMkOyV8RKrUZzEhWVCeVypZfZLlkV
+uLM2q4MevKAUMXYIJFWkvWmAdlex200X/rC03jqFCBC4FNy3weooLRVzF0dA3DD
Kyp/5Qa0uQoULBJWa1gGN7YX+vq/OUAVqt/dHVPVr4j42AfYNjtGiPesobn7dX4h
a4VFT3y64IsjkwL6Q3J+Yjy5NnCOjBsi1nd0xoOUCVab0vDWabMGbokkZS8nwImk
25ts4nh0z57g0zpwV27pEKilqPBf/dXzei2W374a6V1XZ1yCf193C1T3ryqlv+1e
rH+eP4iz9OUKD3IzgIpnGl5V9ZapODMBuH2uUTc4VCqXEzzRqbdaP2M5obdUNrtF
7RNILQn8RBg3Zb7/Kuri27xpmndzIS/w3CdiIfEqwJX1TMsVUdzQZfPnH6pzC+4a
7C8Ao9tdjiNJwNjyp6hlPZdXVnquqMOINZJjM7ZGeugTAAzp0GKyZwdEDf5fThmy
Ef6SI5i4hxRSV0+wv/5Z/bMYUMgedfbgXFtLy6tmoeO7g+k4IJtTnnHhVmkmLP8c
EkFQJPMCx5OnTk9RS0iOFW5IduddNuP6hl6IgfzGxlXFywwpuIr47DNI7YXd2Y+o
wge/pLse9jiS7Oy4+U6twXrbQte5uOIojpKDh3Adt4HIcRe0O8uljpgCN0pGQlsK
pvkKWlTqBDSabnP30euCMN5vox/3B1n9bzbJKgy4ZqRG+BE5goHZQ1kigQIVa7nb
VZrc8j1YXmWfiso16ERhExA1a+V26UHaFxtnZmA/J08XaO2Nz2dEnFFWUFYKpb8b
VICzrVnQs6fBzz96OrCJQJd2Qx6qQ5QC6o/hkeTfaYeM/ofUmrJXvDDDpU/6ktlM
A7qq0XMPiZPxP5mM8nHKlSoCUpcF8Rh6o8zgY3qeN5dYWXUz3nq4gTRl6dYOWn8c
+CtINmO1yVmydmCiztr3lfBkjQuF+UiiP2LUKLTxLV/6mYCtzuEpKhU9zGaOfuAX
EVYirIKvZibWvnc17a89XE7RW1LpWbiOLHYGb3/qUf/dlfpv7vrvbYxVdckOSSCk
gBeMl7pCt4tTuC+8jONJfqxr9EHy7O8UDqvFECvE3Uom/IoJVUxMGyMXmbapqJi5
jEnoMEB6KKvs0onCkqPVPRtXz/m7AVhetIx4b9iWLMHsaoeK0vcJol15/iBg5EEr
3NQp0kl1WtyJsypLblCl51P2xb2RyT0ruRE/em6rGXaAp9AoCBU7HXm59Reo+iZj
lxTHp/61AlmOuxyq4dScpURQDDa3C2SDhfTsq+cg/Gojy+lqiF7mO7xqqbTdom3L
hBF5/wUmxZlehFzVfe5cLxqj//RYbX/5io85AKNas1N5RMDr90xXqOKJ06cx1pGj
4nIsuI0E4CnDivdBEkqrE1fWn7Dp0IC6egJ8i4g8p+il/4DlYw886/uvggQjrRXB
0PbruwIswNK6GZdXjYwfAKlUlwGMw/a80c4+EEe2OmaNf/ydcFXbbSLgOcYW9xr+
p3iAcEppSgdPVNvEFaVschWlsFJ+MJV2r+smoa9JNQB93oXZlXTn/q2FbQWpF0X1
XBxjbyks6K7r8dSWeOOGwdLOi+mwEjMrEE6U9IkfHPzsU7MJVFxaggeIgO6yLmMU
YSjgXgLBcYu7oJf4t3777VWG3iZTZqYBjDFhuUcOyF1GS4kfQVyd2vmZ9Qca3L2Z
lVx8knTjvBrgJ8ttTWn6UtXynY/rbj2ZZkyGBtir6tbftF7z1WgB1kFQ4qCxJBC0
pKaAPIhQT+tCVVx7ksGkg3+cB5IzRKGLzZNPw/kgO8vaSzr1Xi/Z1ehcS1jPSX6u
FU2pCT50g76klLJXQbexiDmz9Wm40r+DXu+YZ/AYTaROoY+GMYLfsjyouHJow9oN
NcOfEuXfP71LxFMdvw0zp3H8G+iFb3J9sy7XuiqQlb4i/+pBYW6FLJALdXCU3FtI
/sLB2Al3KHNFz6Fkmr6LyXirqBZZckORlb8mWDVvnB4TToQej3gpGSuWkEPySa6W
jv7r5n244FL/qT0x2r1zX5Y6B8lnPfsq0JlwE0bQeV0pplrnZCUU4hLfiV6py5fm
V19Jx97YGE+7WmFHEK1zLmXfAnZsErVAUQI9CjMh0HAq2PLma20//ZddUmS7CgTh
crw5jUpReNGEpRNIlfBzyyfNgzfOKkc7CPFm3d0bshja3Wq7QBTStmfQnjLU06bk
EwCWQTQY0pwgAKO6tiuuUsFkehejNCRCpcLak6EHneQ63oOq/9AiMrte4KoGpLG3
5vSm4sS3EfrGFREiDvCFJd6l4gINhRBZ6KsGgmdhzsVVbS0fx1a/f/y1Y53SIXI3
wy0Nj8ACdZQdmFU+Y6SEOmxr9OgRcJGZ/lsrL5IhMK4OMEcGRWRMFZbMwyNMI7ml
rD/w1htAaJFAVEEb/gwgEHNyItBgVR7N+3lbIuPa9HuE/uaME8620LY4mflWI5VP
8+Z1A6MeEciEPOUaRUJs96aAA6fWW6zPACQ20X/vHF+vm1lw+zY6hKvyy0DByoJg
fm/ju1rWgYSlanChclQ4pJlfCz3kRnZcRC+OzQsR7x0NRwvgHG/jr64zTe+WbRjM
AnS6qim+Q4TeS6ExWv01yUJfThCSUqXYe4SsxipG9GX/NyzoPtN+2bzfGc4XGbL5
4CegGtb9VpE/RECz8CnAtrKL7Rk6KRlIqYdThNKP6MNEsewWswr0J+CWbbreqN5J
8Soey/MuvGXx0pb6SmXhIdrsyOYk5RzICFcjeScoDFiaBiruWcIW7um5RUP23+Cr
GrYjGDL8kc4lhML/TFGpEHyAZHfC8LfUmzrawLv6Q4PDjuUnotllviOpyC+aihGa
238Ttn9/eV8cZfHeuw3kBaz/IZJR55R6grS1qlN6Bb5ScYzaxFCTIQCM1RHHLNER
0SyugdbjmL8D1zyqAStgTBTPEi9/ippca3jUxOc3T5jiUP5+QAAoqU6ZtH3tI0rL
m/sKC6Rnj1VZ6q/alU5XiRfszlMtcnFzwAcAf2srZsaXSJdgzGP/HDfPhlb14Cx8
knxpfEA9AuMTNCwLE9aDc6ZhEXcjnC4m5VH+v1FFHqW9Bm/6fyqBh2/h3Vdbkcma
0dANYo+Do8bXAXQbnobQ3CmfHPC/6wQrvzk0Vm+q2YBWJuDu81GmAS8jQA6I147j
g1s4tDUg80F6b3QFdVBotQK7RgrHHJR3cd1OravxKtCbKrjfZninZDCfK27O8sFt
9C72K4zavZOcIV7ZFX2hUXQFcZcV68PXGDRN+nMelpeDQpvXVTFsm/e6O+jEdUJj
WbR6k1AiiP4qOxJkataxdG8fL9qLDMmofEY7XAdzEpyzm1w0hDuM3njz4Nkebh98
Q3i4FQ2cjkYeYNEa5ol6Kr2Y8BRMSwnBCzAkMEp2IQJ//HktFbMOqW+0zWVJvtho
LNZKIcpwP0IJUzhAFDqfe7/n26DHy2+ZONOUOnCDkXYbYLmL5O28iRzM5uSyI88M
RamquXoyNr0LB4t8bKpJeeZYv079gPYJ9e3MTeRNIbEwcCJVfIlYz74u6Eb+25Fc
wJw4cPgra1s/jZG8sXZiIO1CCdBDe/RDy+XgZ6gVCeuEn66iUZomayBG5Hd3vDIq
NKeEcxfJfwZb+ZiVEgO8X4Zv9/uBnkFEF/vMGEuWfJcMPXr7cEEOeCb8f+qeGlnq
NSO6wyJYKZAvKQ6h+6784COasQt1WozhULf7dH4/oqSnNbEIucxfm9lUUogfGZWq
FD/lnRBCRFvOZeoV6UePHX0EQjsq2BOcDX8LdXwvTUcQ6epzFesGmhOgx7HFrBN5
kK9u3puqcaqi6+cjFK14u3EUbbekdpjFQMLDb1qTJAPBGhmnUvA+4q9UknRocXZx
71pK6IZSHUKuMlUGgsUHYB+ZVxoWZzImuyFpDh1wPx6syCF5tfevdAclvnBNYEBt
AUKKui95xtvoINbiuKb3OjsWafFj4MnWOcJgmNA4bNRHltFfWvKE+1MRhXKWqKxn
SgogSKehZQPZEZNGg9gQyw9GR92gfD/t8fq2Tocb3CFNDKEp37dfqNDtyvSSzBva
/sYRiXNpClEO8Y1wJUkypCYGC0KQ7b1GG2P76yJapQcp02tWZIjVfDhqNQ74bgRB
8obpmql+64K0cYpAqrTPu/9jcsce42XBHmGUnIzfQL0cWyxZd+NLWtzclCU1TGRI
oKlUrnPjLVKoRudHJlP8fG4Ot1Yd/2i69YqfZWgl2oVOkpbgKjsQhp4ToV8zUJCD
zQm2nmNmU5R9Pe+FwhjivR4qu/fvHjMtpUapcQQ0WuQ+/mkp2sEtNECou74fQp3Q
eL5gELN/xyXtcLlDp/aLK6lqLEf+lFesD2MwlzZg4kKe3ZvHiv9Z7+1aiqkGwIKJ
E/mLg6FJ89McIIuIaIWPPr6E9MP5SfFXPuZT/D7/2vD8pYFCbuAMhhoT2sOZPgZK
ILS8jkFZrR208/LOWktRgt6AF+tu2VucT20LGsKuta0ZzxsZ2me+evXH8efbf6be
/VFisQ6MIlGVzeoJAKwaY/sYHo8yqklrW1JzmK60x7c3+F6S7gasw/gH/n2ep5aW
8E9FMSW/+/1XPewX5nKflmugKp04CjhYBH0tejT7K10+CfrxRXFgjTZq2awuQ4EO
nzjvBek4KIrbguQ/jQ8wE4a61/B8erq6MZsZwwCJKDIBY61DQvQ5StXowW0t/CAd
ODcY5J7HqeFcP3WkOCVh4z/vJepeYsw19U7xF8NOwFmIHgjs8VemDmp1y3uINYS1
ksFl8jZJNzC4pC5/8e96aAHFTZB8J1STuScJkihXHB/MGfHcfoure6H7bekEqK6j
AElF3Z9/AZ/vtBYmjWI9qt5RNRXxftBK2uuTRGKvLtTppGq5w5HIaAbpCNU+0Rle
klEUbDGRju8bUEYciVzuqAIrzT5k5MOGHxlhwnCjXbpsiIPxvyFy6W9zwvCo5GQ1
Iq6QcLdVfKSvC4Sbz5m1nXM8piaxblEI/DzzfDJ+WR0yhS8+Be+qA9iC4/MIHd1o
FjcyXa2CYBS4f9mvalHgPmESn4Potb52azW/0/Ws8E7KObNhK+7glKh6V3dwNx+B
SGSteEF1FiftN6hOQpwEZ3L/HxOKFL++d1WziqKsyIIZ1cJGR/l8iUhVCtiywFty
8cCzOWyCQLIbMBVNB/rVaoPB0qTh+Wly7dJ+KOZWiGy/bSoPQ3lP0tTyAAPondM5
ByEmNm0G5yQmeciPKOeD2S8FNGDVdX2Y9thNIwZNAIxeEBHBeXSDaxX5NaJQpdT/
ktSfaWfpIB1rVR3sacJhz6XAoAFrkC3x0ABgAyIpBKwpa5SAy+p0mCkFmA/Sh3Xq
yDb3mD04v+XN8OqaeUxYUzJOTIgr9ypbgVl7vUQZNMJ0YqCe9NMsaMlx9Fl0mW/u
y6CzbnUUH85E0GogXXlqrsY5wP9tEd2cM6twPIGvfTcN3+bBqMDf0AR+prUiiniT
AhTjb0gApS5sdLnVisPiQTH1pLSBpNuuz2yJz69H2nA83thAUfHiFwcQBz9TDwD/
V4CbXsoZnmdU84Ap5VFK3IOOg5tP2pJ8tPs0mIhqbFNKkiABhMFqnBm+ghG291mo
QL/VpmJYBRSZuUU9PqheKWjRYCwuXqsZslGXCPS9TYZhHK5xLvhWdMmN+BVJvJkQ
Xdy3EfDs8OUYswtGCSDS2k6dGw1DpvYGlMWW5DHFIR3o5UJZjNJvQXZUsVSJewBH
3uUoJ9WwcwnMwjzb3q3GKIseCT08V/ApdElq1D3BlgjFoA+a3ss4YRZTyBg9uRZK
iIup26nIpVhdGzAwLmaYQ0vIvOlkEobXrlj5+O3GBaD/UvtmtI67BVXeOEnQoxtF
pgTedC9a1JqxAhUpxxJAAMXunAuBBR+aHqXoyHD0c410pi4zXAQ1NkC2ieyXG1Rn
he2Q3gPG7qHWWYxLdOCqmvNf0o03qdQbR+hv87/uW8csfq7UpFHrczc+2PxbCAGc
WvDq0Qc5hJXxZlzVBTUmSO85VfY5bHThzSs1Z/XwO9/Q5TTy7MOUxSQ1dBmpR8jz
msoG0xuubNlpnVmWMTSLI2ePGqLMOdtabswGvQqvEpDFCTJuj49osdEbxf1jP3GW
5RMEWSnTrzcJVrCzYhu+i+wRf2pNKVRQEnxWfAiX2hDGO7v+NrqF7ajN5X05l5I7
AvXiVuBg8JRlZJ0cW0hIaMoay481a/Y1elu//sIJT8BR6dnd9tgNxLQJuigEnO0Q
JScsLD/gMtETgT5O2ONTbFMrt1erv4QMgnSUKR5znEo10b2qQ2EyE9BAt42103WU
Ma/1FDDD3NXCoKkoqg4oGxbHnrEGj3aylJejmji4f+skfOPGwd4RuIu91sHGro33
RhTssRSLan0eOVaJgLET8Igv6XmATxcoxvSxQodtszSkylxgeJtC6f8GUN2j/i3J
ecSGnV+LHiRDY4q51QI1aM2ZPosSc2uXD2ZZsXZT637QPwJWVdt8GhPK+i/jKC7k
80JacJG3KLDupH1F3lRsXwxafLldmRwuLX+qg8wRPrcc/oblsIDY2SqEddFj8m2k
MP4/kq0RZGTUFJpJLv9IRCwqg2oJ98lGyjdk9aipilxpncZ3PCcfFpCAl4LzgvN4
+SoI2S7HUWyRTdMycYCuyQwslSVfHxmh5FntoCEVa5Wn9mJb2DzbRGlseaocM+bg
aecqvILKsYwqZJvXXk7Kv0Z7whCPymCpPiLdXbZO/fuurkoWW7/9Id4N/EGVB6BP
7zozGyZEk2mKJMcJijz6ZIcIM/D8b0kztroA0NIA/MPlM405hbukLI7z/FKOcKBs
unuRn/WLDRU32OislRBeudzYLoZPdgY9JJ7h4o8dD4E2GrNcr7pEc/8ncYq1Olba
sNKBnREzAJDoHm7X6g6vmi9ZNvlsrMqH67+UJHFJZlUYjqRQZjKmcMEnk+1h6dTz
aNKnfb+QxypvxEG88t7uiZ3TM2AQGwqJbs0ZICA2wdZN1rEmJQUv6Gs7RyivGL/H
+kT2DwWyxbrGkolgMsyhHZXdtykJLLMvRAAHUpPUAVtHDmVHY8ChkUdwBgHRNL8Z
1Am8stRhY5Zd3uuCE+BGMN1dbfTIENHmkBR2xEXmj8dlP22k+RWtCqvSlB9ovCz8
EaKAlVq2QgSA+1awk+IzL4NE4eQtPFZTN24QD747GKI2MZHSlADwiHxRjuWk6PAs
yRRxb81ZK7LL0y14tEebFKcaKmUH/MDggXiDTp0jAvMLcr84FXuLcuvpchBiyo3j
EoUHlaK+rJU/HoHHkCh64N6UtXWMzqbk6/joSxe/j4IlzivM2NTzTLrIgwUwqi7p
yY/nd+cPiosaJCDesxMVO8zF5hceB3Xir93UNpc0tr/+YVpLOTNQhzmOKFzPl5C6
L1CeUJwegsAW/ONNpByS8M+zTuNmJbwVIPnpo5YYACyh5cCYfw5+LdPw3mCB1Evm
t3N/cse51JUEU3psmZb0V9bJAIqYgvbKUzpa8rvSRaHpmPnE7UumHGGtq2ejA9I/
Wy5MnQbusxJkzhnHfxfNZp2eZsDZ7ZLvIJwDTR1iBNrVb3e1joqzc3Bhon9pYr5+
L09qnBpkxRo1/nIiMtyRR01Iz5Cyj1ElKyrbOLDRVDr4FLb7kASOy1BtOPpq9rtX
Zfsv607F7TsU2Wa3FEtvHpQpqEtv+otlGB1veMFLC40qsYd94qF7q4UwqJN+SR0Y
Q6xtI+knGi84PmUHQB4YzkLjdGDROWaBNJL88c3XqKSZBA++7s1syY4mgdhRIrvn
nv9+8t+i5Mng3QUCJ7hzSr1mcVTizIbgeymiFmstfVR/qN7SIZGLYbMwybJb+1ar
Gg8uEtrGkDe0j46skBLCS+RxV8xSPxRRplKHueU5jAlqi5G+n7VIM+b7i8iV9FYV
/qqryJ0kzybDLus419+mMACCU5oCXEuY6tzNtpXcPcNdBr2x79lUK59pV/5lnBl/
Vy2w7lVt1iT9077FUcJ5ZK51BUFEr1ke0L7mos7/QteA2ilHVtyd/oV2KrftV2VB
DhhUHl1CuxEZ/1cxBv3JAUwX/GhLxdL/RdJlsu81jtqbvgpQjKTKySLUKhTADUrl
+/SAvOpaACXf8K3xhn42qXSWwnkBuJzHqpOrxFjHHoGdksQrhmPw6rnfUlm4jm2U
PuaCAS3+RisimgREvFkO74ujID/S6ZocM5xBsVBHuW+AX0KfOfOeX5sDPJr+cxyX
6tIjkYp67a5s/3R/kk4+ZMWTykpXDFN3BgWoOazFSCEF5MlkzlsWK4ExdeZ6bYsK
Eq8l3Olrm/PD3HS6KzRApFy8TFsVJXcLUbHJqbEcQPuWMgHlk/yUyr+Cc45oS82T
kntV7vepY1sROc/KPa/BoxrPhFWEQLQA2MGN+WDXzefmyImoAqpAVzpdQqer8tV6
ogEZhWJ1slvmH+OTJJNkI7o683xjfoHG3hTfy/2Ic8nk+7VDZyGTT08O0YjAV0ts
G3ky+WFxU8nlHGAO5meKtITzNTAtMxGg+s780wKrYrqZr4+KR2h0elHQ0XSJlND+
t6A/3VkZzxmq7RJjrgFFqJw06oWC9y3xiZPuITPfsR80tyWhJ+vgKPwx7eXYrJuL
J2WK9OVatbg9UFQZ7YaOuIKHq+3C1AbKGKK5NwcXzh5jHpTBq8COg1dBbxvOIdEO
Lr05cFo4YpMEC5hhJXK9xhYi7lTjoV8vVJNwi0JVKXXzeY2lS2xSmtVpeX1NGjSW
aw1UR74vGqSerfANato4Yw8GcogjPs0okQRziVj00OOxw6JY0C34S0SaqYbhwazH
+dSqccXWSH8dTWTPkFoJAFEzP4cjy9JTXyZMMiUzQmMUElKXuwn/s1Wne96FPRDm
3bL6ZvtwSc9wycS3NXlrrJmq1qx3p7N1NyQCVpt5VZ9XtgaIOmTwAcwBF25VUwQB
KlL7BSuqD0L8lQ8h8znjfbkV2IIR9F+wlmf0NYX+kAzHkpg248L1qFrJ2wqxTNPx
rUMQoxHzkHrNMqd4WJmqFBB81mMC8TC1oI88HFLQQworJ/tlffqJyv8L5eR07rDZ
Y5O8SemBJZSzN/Hhuco7rjnZj692sbOsqO1j1XbF85spUbpIu9A430k7uSJx1/ZA
9ECckgAd5p8wlksZCwXoB8qL0W7s70xhJUR974EIwd9HEHMsKW4Go4HT1AMGKDz0
nk4eTn7kCoqjux2AOSJJ6AJAotiRLpAzMEiX58tj/Zfgu3qp8I3QPUNZKyxGhde/
A5nCOJuAYs4XaszXcHZdZuKJO7ISq2juZ2DEVt9EHuuzuk6kQdKUzubJfORojNEw
zXH3m6My3kbSzB77HDU2wApBhvVlJak+Hp69UIvF2mKHEVRS2NHsNCSkwyRQJ0k0
LDNrduFWEqSRjMQ7mPyX2T6JVuMiTv724Hw/SNKTQzdkxtCiY/qxTDBbuX2x64i2
C18fWKbxZfN5X8Q9wrqV2nZTbVoLNKrefToBAZuoJgrOm28U6bUn1ShpfnM9d04k
ao/WJBgtye0UXcMrtthS5V3ayu68M7hNwFpvQtznWwK7u+fEA55pfvnkzwXfpImF
GgWU/hHX0q1T4dlcc5qoWd7GhoOyplxY1uoBSbJnvALK9b7PZVtugbGYh3MhlmhS
9kfhHofy+8KlfciQ72azYl9c4iU5g8ir7AgpWgPm43mn6qXoDUE7dedUOpFxzeiO
XtLeu6u/0pRtb6YaX9BDoCp1SRlXs0AS4RKlPxVm0I1pLB4TDAjF+WHmGiro4EnN
Mf32P81V31+h00ewnK3Cfh51Rk20x2oxuowZOUXopy+M2G+YvHTS+/eGHFre4TI0
SdjDnajDMGSzFnBL7Ul29Lqs1hl9MDYGma1gbzeJQ4HCZVWz2ytXkTiaxiUBEJGa
+XYT4WGLoy3rXk/by3XSKsrymLiPsKgOj0gLRVGtT8P2Z1ujorXybIbm1m0U8IQK
4SnaWCapppwbSH9pmfSthR73FMKTIiMfvhqNmKZXhueDkV181tGTCy0uGpElrgbF
4Tp4zTMxP0oMHZpP2sL3ULN1wJUr+/ku1J6563nSejjKddt2jKXVSbOdu394XECN
OyyPpxRyhkbuik+SbN3NPhaZdeRZ7hAzvsExUsnp+CuRy7msE0QlZtfJPU41nttu
BCkr0vz82lVMNqM8/Ky7uVE8SKEJJF/N5G80cwGy9Ocb6wc+lqUsZGWEfjivXzkg
QTiUnvh5rMdjQ54yJf6Hzl6XzImTj3i3DY8LBliakRft300NrFHpAqSY+WAmDfxq
DSsUs2XQRFpATKJorJ/QxQlB4Zh8KjObUY2867+gnUIFCDBNeBVNXbz/Tmok7c/P
+UcvKaD7qDzswYzXV1/bHeKGMpQlA2VRAXUofRybReM5mAH2xIcyrDK16nB8M8t6
FuMlgCWxD1Av9dNOtgpsirMVojj/u7FjzBl44a65ZZfUrjNOJ0p0HvWJTGDqsiwn
j+2DOpr6qWN2xn37Mby6U0vn0fZFOBSXieSGY6awkGQznyy2qcubBECzsru0Ib+s
YhbmjX4oZ+6PM3HMaRdryBW4OBDrG/ErNI+BETjjr1DURgvu9AVBT1gOQ9pQ5Ov0
i+TCY5q5Z29Of66ywjwswzcoLABx8Zgu63BgRBHD8QUETaErl1ebUFgKoGruKU1O
c1JdKIAy9N5T54bW3TglhpDpD0wi3RDM5mVGs57HxzaAoosDI1IrV79t/NwXQU9+
CI+P7XqCEfEjK0hI6L81ckQh1UQn4iROVEFqtDmfwGHlBVjVMTvuV8cPp0DFqZkz
SW5KNXbrMH7pV54DsinFb5UcxhSahpMY0YfLMVW7JA6lRS6q6i9wXlFhww257R8i
xQAgllLXF8BYHQk6sq/t0P7N6/BM8DQIo5YNdUpI4O/JwB6ZmbfumiCRsJgCCA6k
n8ihxjqiZoi5lxa5E1oyxGLww5mVbiNEyrfYjRmoO00GWpvf+JEKmA7iFYE2hW8x
kIAjNa1R+tUvNeN9wQCMeSAykk97K+Xh0L1n5i4gACn4+YNf34XAq3SXeoWE6BU2
45JrEsdzfmZRb/xBCpXlBDKnu+vQSsNu4igirmpUZbwRJ/X7GYcpx7SuLq0rHxHe
vSgrIZdnEn17NBqFQdsvDbCaVrYY8AveAhbn+XMiw5QZSeFd1qpSMuAR9b3w+K6D
VqhAPaquh+8j2XW/YY4UrK2ZmBtc1lqPJTgxTQ+zQ+r8z1L3byOanrsZ1yNQ/I8r
qVxjswg3JOrwdDnRiY4z7ZSDcM82Tmbbj7MD8oPMXqauvoavW+eECoYTwAISdpQ3
+eBjOK4Fdr48JJ2w3brPgg/+Op5wyDcZEfY/HROeZ/vHL867l6XBIfbxWde1Bire
rOCttYP6OhGBAaxXKjbi1nGsDfPLy+F9Oh2YdjgSRXQh1aPx6lrkENVgfdVxeYAQ
TWKuTpFEO12gUub8cmPzT/dOzMZrGnSPWxGspPVwB50aDqlN906p6qSvUZVii32N
m2mAjTDKL0a7ePqIYkxg27wGrPnM8Y58IzGLRJK/+d7QuuQ+FaAI3WoMGRkoLSYP
zENojk2vqRE4SxTbPYTHQkacdBnTSMazhP2VCBaju/o+4RfuG3JvywzsP9EdDYCM
598GUvNUHInkhXgbSI8ITnOBZxaF1P0O8d/yLb1Q0EnsMMDXoIDROwR4lc5aYLxj
9cczD9bx3yPGSzeYIW3j2LuxCFMgIzEibuEnYtPgvloFUJWCiH+YE+vn6kXPuXsU
QgVcb0xRamFEBfF/H51PrFCxYaSzqpLkta/oG15KI8BvE7qZe6dI1fn4oiVT7FRv
cH9AtPzlzFAl9PyYNTiCTrCCB8xbT7WYNHgoTEWvR06sPfZZiBkZlGxhWVmk4eq5
9a4h0t+23A/eLfizdYQX9oWKx1lS3d75S8+1X7PpyTT5Rl7QzJbNIrbAFDZ9nSpD
E/OFvSKDRzk0ihlcR8zqBu05HwRhPrS1nOm4IdTJO2avt00mj/PXLI6EpCM9dlXO
Wpb903V7FvAlEo2pzq86cKuXooiTrxQAIxaOZk5gWkV4e0gJNJsdjGV4DG5v0lTA
IEMo4yXaae1BnxF7FZwigoxC6947GZlN1jcfeNbwpGEIJVEO59FExqGDPLYSCP7Z
yRjguHtmwXgfmyT26gDxgn9C/wss6nApSii2yRnZKQnBKly0pcxLNDibvckjlabm
69PtFWLADjucA4s+PZxTv77ETSF5xAm4ndIVQ66zvs+wq+YTukPKvA9q8i30G+TI
5dc3JQ4AFLgIlzE4AT+Q3vaRxKUo9BLtbdNjM8n6oLZl/ddyDSbBA2cfA6e32S5s
5j+OYDgg7YjlOiLnSfgRpnjp6c4PRh1bbifQ5jv9TAmDyw21y/xw7qLYo/OTujwS
1Ou3u/zK8dFRQPNVjr6q8y9EWuHoW6kkX2QdBL1OBN4BWRCjhfcBSaYvUJUJEQVO
ESKtflrF6xP8OwfNIPE3UvptznXO/tACzc2mUGMh16CWV3vWI0CgDH4WkITmrkFP
iyGt06mufXXhkTj4uY6Qnv2UMBT3XLAI8Zj6i3IoC0UvJY886UqiJQz3fw4zVFYJ
RftiET57rnpPh4QXroPxiSg/ZPgtUjZwuUEMMXj6cii4Q9rMPBk4I8XpmsomPQsu
r95eYo1vXQbejQgBJ9rQ1ASdn82oUyM0QTFEfWJRqXm8vOMOB242/n4sDdfxnbYn
LgABTn+wfS8XtirqC4WO7W40Oz5MNC1oI7b33FnMtiFRfnmmAObBJj83XKMo97Zl
QdVjmiDBDzH+pLQvdcQUhhO+7CdIOIyx/ZS8fY66rWn8Kd6OyNEtkx6MD+eVR6hn
Q73pRUHz9EGzNNKZWBTKUJcnivdoG/wyXXiYORrZDhfsyJB1SbGUOmyu4yzz+FLX
t5htsiHemOqI3Gmjz0CBs2WxGZ47nQJlDNUulAKlF6XSZfAjxn5tbk7TUsS73aD/
Mc6OtlHtBu7E8NwaoKgH6cG0sytbq9uA+X/Hn85m8rcgPGZC8+RZiZv6x/V8oST/
wLq3WjDKAxETGMq94Wa/hJ4N5vt5Wsk8RtjOD7/RMfwU1KCiRSVqvAx32QbOhOZQ
p7kio8lxXI2yxtzSDTWyOEGB1AROg4FjqxelzwDUojKxt/7+Pt6j2zb/2z9Jwc/R
QYwoofX57oeOfGiieqrdE8BYCmBqaxKwfNHxREcXBOzy3Je40ewcyqZNG+HPI73S
z89NyKgAx+yKmwd60TslneaOqCkLIXFEitKUlWMvkYHPRRR+fWC/1kkoWl/l/l/d
qjg5zAM3KtoF6rP+9HEdZlglhqV/Js6U/MGXiiu3DqfoCJGroEnswHarVICF+Ly3
mtqJdYLprWrOLx2s7jYy2VxnHq/FeRY2mrp6E/cqCTvdoF4Os/0PZhEWNrnc2FfE
qpGE35Ho/lavQJFWW3qoHFWnvpFtytaguxy4SlorBHQbinA3YLxCL5t3chrPkneD
5EBP6pdQJ+oBCjeOBGvl8b/sdZy2ePPpOzNKfwlfROwbpbNzsjY/dyl/KEk/S6fp
VMdSzc9BXWGUnxE0/Y2vBeISL0o8oXul7FsNATg9Hkc4Jw6r7/BDK2M+1W0QKHMz
4dXfy2DLie8iuwLJIR4qmoTISDdxiVgroBNu5efJEVj4btzxVH5azvPi3BV92ILt
WkPKJ0gxTcB2kOefIVKeiR/N/m3WqRHVoQ/AkNJKtEecLM6PmTsatwjOoKuDSYVf
y9HSIZOQurOMOW+dARz9jMYYzBqfB+6/g0laGdXiuGxU0A6a+dSbHneM/cLzqYcF
+TvXe072EzHHasmMdaU5m7D4M9tDJqUloHb/qMc9/ApWIZwUw5iP4x8nwUy6Mldi
z/Nc66fTBvKrNk07NbtE69PimDeDV1a4bw3kkaR42kKmNWrKaRPKvVyoYiGQVcX5
nbh4BfM5VdvwYkRU/SLjaKQSYJyfmoSMpwENCflbVD3yRFuQ8+fuZhdHP1DBuoeD
dHXazBmlvuDTC4qoIrmwu01GUiAVbsLgFYhG4mpip7VizfDOE/b6NNaK2YTn5Uqy
zQmjGLtTWJuKomDhFP5FoKGD6z8BVs4K04ov2m8RrCOOouxn+/kaMbD4PW9B+JpT
xl103qVxQiRIMfpDwvnSKVqX8wHFAVd9VfxxWICvvuUHBhVD1MTFEKtrX8onqbsu
riRFDuIWKaOMJji4CE6mGwaA1bv2IOs5TjIUchKk3U0Cj6Mk+VDrOF1/y1SiiaRn
EK//d3TYf9gvFrzdb2kmDVlUXJXdtIU3pOVtwTYwdM3AcbG6OAnTfMyBMmEm2pTM
vOJPv1DzA6auAhCeNXZABtEkX/bI+k4qoLX7rL6kvSvojK8w0+qenktY9rKOKTxQ
cN+LZC2ETJwwgqHt6PenhgTKNQOyKlyuSYHfUiE0aHwIiUpoY+GW6wAOqFBCLPJ+
8dRdQfKprqpkx2fSzeWoJTcKxBiOY4K2jUWbdkyEsqbUBCr/Dfui7YTRjpqWJuI1
KP4JZEz+1yGT25AMWoTpBA/oFw8OVh9KBZMhtUHJonqGP17WjKckuzLRSbm7ZEhk
tmOnPsufQesSHb0y/SjJAFFueZbWILCGf3eLl3c813FokskgG+hrhHTFbIimIaan
JHKhWjD4TVfqWyPtM1AITBNNfarkfXe2dzvUAv6sJpEXNNo+WBOPhkHO0q8iWWYm
wHAP6Dvmx/TmI5RJtxHifta9lb45RAA23ysX15vhqqzep62cP2GEjcupAIUAsXpN
JCu4B9WNbEt4RQkE2fBI/Dx1FN7c8smVSkDCApNYLUkUUI3Zr4JNrQg5V/JwGCTG
sGPuSytKdUeKQXD3ETsuJSGcGnUfe5nOmM30ZjYJVb1QxVmOcD9e3zBdwIFUhnyo
zm97HZf6j7D8qfpctyg7sVe0OtBP9kXqpg3YGJFDkfBiKSje2VrfgoyDJNaHXvcZ
5VRAAF+a99VjbXuxXkga/fpT9uO+kjhIiw1mKZrsu/ZI1ktX+zvv7O8cZLaR61TR
kOsTy4A1kA6O6JGu2JMftUQyAEtPGNieADTZ7vbVw2r0FfJjbz/7qy5+aAQc8BFT
bpXFFASvj0HGGOQ4XMyk77sZYLj/x26bCQcQNFdrwR4aY1fUq/fCyx7DCVVrmmeN
UFzI8aDj2qQXUgz6qh33pAL22L90OhSELUQoOeo7XRXT3cqNZZjCfNjeI6EtxJxv
wtURF3PpszK7KJsyn1fPPD3ABAVp5OU3xADYBl+8QJ7AMGdzkZBYrdiTYZsYfd1d
NeEFkNH61jtAibyaRAOdsqXr1hRT/QTanbntRTwdAnTfsdbDoBZJNQDnTpjOF+/T
/YDi3Ngl43BhIOVHL5lZ6vPX9pCEZMBpu+f4fO5SaWqDTnckCEO54xHPhTO3WVPH
GX63mx+TVHID1kpRRUH5PcQ5Y3dfRXFtdr2A2TXLNIUyFThoMzyKdkl1/C8R1w98
RbActXirMhyzOwLP7KlLXw79Kq1SjfwuOK1jmIXsnGXWlvVsrUAAGvcMTp+a/Hq1
BZJPUmP/kcsXby85/3Dhz2epy3CC31qHoHLWpFkgXlRvFM4yDZbrDGoVCKU4djRx
vAKheqaDb+WABnrxR7fx0L+mAwSa/KjpQ+Y9GvOOQdfMU5SxRBVBvWOWfOuoODJd
/OEDx5j85F0hzkfqbhRfMfcqSXJQd3Mb+Ar4dKE9CHobAzBSBG2gcnWQj/rhQO4X
atYaY1mIreOWiN3y9h42eNr6ACcDcWcimHOMwHjtjmG7dd78eOSXizymqkNE66DE
Zn5UWWlTZ/u0cdJQOmejwYqd6/6xHHl1mxRISc9VHFLIcRtBl4AwmF0L+aRyKnUK
dEG1HzrUXJ1MjVUi0/OfHFvQm73DtEbYFHdKgPp+xFlvtXssXIVTRN0uuH6rEEyI
vPLoGEYRmRuYjrxJds5VObC40Hs/0z0X3HGnLOGmAiEnDnEVriUVMXok/uFIKG2W
qu7fBxkjN7qT8hDZMRFwgELq5eqAjWHgI18ZARNXu8LPi1UxzUvRPrMIeUQrYlZl
BBycr01iB1mP5EZNsctEGMi7Ow1SMX5kVtHuF4qlEqpgnBwk665KCnXhHBhuySiA
HPA4d4zzdAzlzqL6NpI6jd9h0pd0gCmR9YDcU1VxzVBC5Z0n+XyLmHRGt7IxLjJG
RRuj2UJiGXeb8ZnL1pxFFAYlBOSzEFmHS9DCdcTzOJiwLteJ/8y8lC404wNBBY5+
qUpHI9wa+mGPo2yvNjllRAxpVAkCeUvJxgUoL8d+jUwLDqrqobrxusvJ2V0fbuHW
6mEA4+hti+qdWGtX03XooXs/Z+mGAg6WNWDkQ53w+mfqxMZnoAzHi2TKei9BDsvc
1oZRWNOwPmxFeYj0Gm2gxauqi/4inLDngG/QgzHRZStuBVpfbkQdt2VZUOC3X72g
zFHdFKJlc+4jBubOz9Qk9CjFIptj4zH1PpNR9PD5+ABTKqv0bAgzhYZ348dHoxBI
WMB63uJvpUMEX9wYi7ZsPTgPoJelofYqgDZ9wPeQhzNHmhoZFzmtQv2T03ZFQoiR
ZVopSDoH1fRIUzbYJWQm120uGllsL3UP0e+tAuAaeR3nNyxgWWo0WT0tPgMtjir9
wx9snd2HgZ6z13TQuYHI/rRYHpWhiblKasNGMwNRJdzdrC3ldZvMFod0lS9X7xbz
Ot5e9vVGHfEjOIM8M+1erOfQe2bi7kzrdtTXb2S3SKd5Gk9jTwyoxuD+3KLN3BOF
KMpcgKoINxjylMjf1AfdwEOha+aYzSesmS1I+DRmSrc2w0ksRs79bkrIz7TVvcuj
kToxPcjbKjpY4uzIcgzGSIDmK5t2nUymIBlDc3LiKpoifeZh6/qnxax7SK104sso
nSG/p40HcEn/L3AZbjR8b1t1skuOX0rG6NU8OmedF+nQoJLOQMSo/S/Hq54uyaLn
6xaGjG4Yu9LDNAWfPF6aab1qCK40sJfqCJG27t5SraFN0Nq2vbyYb6s+4HUoguRV
osiy4u5YbjQuiz8MxXu/lPHGHLP8WOHmgastWfFXqpXUOLBV7upCRt/AL20NCxoV
W8teSSOEGmeYm9+/RC3V9jfqLcd0T+54tZAdIL80YzJyfJdkE2Yw9Wfl05q0+csw
XIsL1lxOJ3Rmf6wu1e51S4bhv69BcD4ZKvAoDBclAd/c02Ygoc/6KME1jSLMQ/Ji
ZF0P90oIioNtYQUj3+iiBSrRWMI/u54amkZl7OOR7Ka8YN5FKzNz68DVtLaJ2iUv
0VNlnf02fDAuA4uMz8W9ghsJvOd/5yc4+nX+NCNeF/kLKI8rPR19reGMF4dCfOVd
ZUyHD0SUHZE01sajOpDKvBEOdJKD+GFbwQSJ77igmHRrkPQdXUtwoEQsyct3lWN7
prlBMOUpdRS9cGP7GDDvFSjegomfpQQsVb44Plil4UMQi73CFu+JLu2aFnjyp4UH
K+5kopEit7I3soXp+lOSvJRMTg2OOpEHT5r11NSp1d1gH95mLghTiqzHuPGP2WBH
lxOysfPlUjzJ69jyMR1JXgA8H4TRyhPN7vHolPd8fmCxQ/SiiE7V2l7JsfqVitX9
rsaIC+2Q7ouW5rTEGO0iwxvh4GTo1nEiTPWiTq9KmHzqMTuNoZzYYxlLvKPc8HxM
jCwVi3TwECezgZa5Us9x007YoqC2XA8mGIeUDaaHe/g27sXQonFL2RedI82oZRzA
PvckuQ72fTM+1fH14RzBpqpxS+FCt1qov+x3AcgNNyrncrtaffd2e3ZMhOBKRmqO
YEnw+1cysb8GpvSZVsV2518e8sVsNRblhBPPK8mvcm20nVs951ifZ0lJ/ZP/a3GU
41GiC1CnSnOOr/4Pv6PjxXF4ubWzlU/UKvO+N71W0Y0tzFPIm0+8izacyMkGafSx
porh665E29S9q3cE5F4XTR6T54zFqYF7/AGLtNg9A8/kWPPz4k77CUR5vxq8j/47
NPwCYxVIaH+oH6dcpIcxbzDY6IhnHFxVx+RFrTrVR9RfVBQpd2YxiLvNEZCbEGWR
kRBrVhQFuPJ0veJEEo0WWJBsMpJAdvrjJh3zjQ3Rs7FjYOdlQYfdVHtVKgAMbMk7
GtCdRT229bkSj8/7dV5yIuxSMWEzvh/ipftJ4GHhcrA/ECMjJZ1pdmzwpxkKZOQe
GuRhLZQg1yBmZ4jX8PtJJjwlZ+6wNvKvBJY9MW2MLNanJ6SbNK0UoNYM8c50sTjf
ViYpvYVGrVp3AbEji+qC9SOGh6P+dy0GSZFlrNxYIItAdmyDBMw+1psIcdI6y7FU
wzNkbk1WPEoik0ATPNgTVmG04in41H1yxWA7o/DlOrMSJFeeCS4+ZPQP/knkMhys
nogPCiLURDd8W+/D4czaU6FimTJ8/aprEyIqm+uu3K3tdKagCvUy7TYu5CyVQSm7
S0UHSrgnxTrtS/ZwlxF30oTRuhSHBDKsgOTbtB4o0ybZ7iFPxcmPS/5ae4t8Rzn/
lYR8rXVRJoRY+azviSNQ9TSYn4qnvlfBRdJd2XI4RuY3PQSo7Bf+fngzMfQJItLL
5ze5cybQsNRvG18ql5Pe+3dJd9M6oEFNbHMH0JvRxj9oOnQl94jjf+HkfcQjMWye
XKv6vPHiow+4RHulBPKgChc1Ogm2NLLmKvccPbzAKtOaDS2e7aBpFHWY5oFdOVM2
pAwktvxt35/iZGc1paY6O+MSZ3bVgpwBKHZTzKs/AMJnNKLMEHpDM7p9aMMKIPqt
AopTrLRBgR2ojqJ1J2x/wZROHu2UIvGESnd/s1yP+3tSvN+f34mXGExwayHvh44w
ax9O7ZMaTaYQFlonsj6UqJ4nqTXG+mMCaIfEuYVklIozTCbTRwUtg+Tu7fHNSjyk
m6ziQY+nUYAW2nHlyhgFPR+ydBjbOWCNgWY2vPH+8kzZM4SlByupSjGzd4/lFOPv
r7PDQ3U1Adnlrz/Wr5IoBEGecWbf5YiG0N4xw3vQpjp0I2CUw229GqifNyxLPHUl
N7C0XzDVy73EP62OvVLpFgnNDkc8SjELNx7pMKqwJg8z5MnLGnmf4QBGyEz9IRby
lYAlPYKCqVeHXhdzp/dSR9y92r8uX92zn2UpaoQXY5FW/vi0vQwlET/QZyT0TsZK
7E6PBuSwo1OLd33/Ue9F/xTYsks1uzRjXJdGcCSBEk0mLs2Z5H3aJKErGdUaJ/4W
IGnVSewmHqyi/7vPcWKty38urgjWiFKjAiZJ8tfikonwh5QAe+z/+hf9vbJcgTdC
SpYI0z64uSXv4gWx4jRFWcYpKUFOiFjvnEtOXQCr5IbJTv3cGF5syAglgbuen0px
EXq1+WBD1vp7jkzxuTyvFqbfeboxgauhW3ngifM0+SwCVCD/HS1UfgNQyfdrxIMZ
Kp8YZo0BlLjO7bWP+JXFhpui8UweGq4L36K0WvNWGIPaswGLmoIe4E21MVHVnzlr
1Cl/fdcFtH468hF6fwT+09eIuqFfaX32JEKIe6atH61YYTY4EOU7i/KsBFhsXK+v
VKFN7ZTSQhc4fZ63q73aUMXmWMbOsMGyIW0GnehMsTYYCdAxjCY6bqkf4NXnKmXQ
bVtklB5ptzUc7jeEts/wcVw+IwE1BioEvUlNKoS2lp2qEtCTWTdcwSD7QRInXkNr
Siwq9hqSxWn1FZmO9DWFxhpRdeQ2qNK2hX4i2hLVRV6xd40sBcOxvjQq090lsOYX
M5NEDj0y238rlCw1hYaqrUzQw9Wtx7AEBKp3LUV4Z1mdtho0myGhRhuIX89MObt5
Homnp2A2gIKuPq+7zgd2W4FSltGJnM1L7G7u34zyRyxyrdpxcHQRlD65afMPSpu+
FSVLQXg0kmJwKHkZCveBT8jAbmJSHtilRqhCOGJz91WhjKJbYtF6xiFrf7ycfOcy
JtkVrP+Z38A9+q8dbAK0zmCia/mRjpwmxNZcwIBwq6qptDssibgO362M7QrFQvJF
WaJVKpyNStQANyZfcQ5OsbyAsarnz4lFfXOzZ5Jh76ARB+D0aOg9baCVKhBKgkcl
G7V5y3OdPrc2C9OqWFq53zl/Qo2Ko12LFTO46XH0I0lhNPanhyBvGKxoijgS5G0p
YPaYyVrDwWY9drIX8Uua8DJKSqVkLCWMLVvGbL3NTnL2enavFG4ReufWyxo4E/+i
2QB8eCv2BjkuKFsifNEkaE2deHpycmi4AXHlMzpFN+4H40WOTTOWyd2eDoXv/8E7
0SJx+KaIDHZQIFVlRtedldMrJebj4d/7DHm1bFYNjkTdHxh7QVgpdY1ovVdVdsNO
6G9XXeqBa9gGfX0VIZNgZsJKOAGOSByncuarLKe31xwmbps0wFRpUU0X3fb/tYbK
boM8bL1vmhmYm6tQ5SoO76hrJrCOwhrscTcvN7F4g/est55RyLQtiEVr9rvfiHST
H12ymJG75nq0hT+RjKrVSXQYcleAtgFs+DqiiRFwpdsMw2W61261q/D8wgbaPRo1
yJXxVJMoN9qlcXsf1hpvsy7p3gYdXmlsRj8QTWPmzEIv0gKzAtXl1kR5+HB6SMYq
6nXWrEPPpQKoRvGc+fsC1hidlflxVWiAPUOZhKcFZaOdctnWVKpUA/CxkHR5XIF+
+giaiRPJG2rxg6GWSGVQvceGfoALEBUGq5Z0/S+GDqtQHY41ZGAA3W8xn3SEGgvj
J5L7pMSMiVauM6NUXAryrdgU7Ohn/HCVYOqjWukjUZP1XjnCePVLZut2Csw023u+
PUBMozjcC9iQzd3dkULYxxInl+QL6O6TV+hA+1781YoloINsHMdbQ9yksR0fVyKc
AONVCff0emhccRhCwHAaNXEkNAqWKCinnYS51FjxvgxwEJ6Q+KSsRW3ByrPTly6l
AK5zsnGLw3Etk8Ddpd6e4Cw2nV+Op/pkj0HJQXK+OC14Jhu8MWv6BhSmZMW/BLRF
39UBkIinX33YCHBQh+5kNFlzQxwSGLAPJ1QADchwrsr1FXLyE6gm79HKf5JjpiKm
b8hhr+8Zv0AMwMzRwF+QT/tZvRKMjEWqlQboPTx2VUZc5yslaJpaIslWtBDztlIL
ZuxepHExR843qyRvdLo4JbnA7BXTA1LiRH/UZINnxENyZqvfEdSUktFEn3pb7rtD
07Tjhpo4FJTDBEYf/QhlDkn9HHcVuwcIlCy+g5ohhCRdaCDSxEBoWBawPIJeLF0I
DXjxVNTo1UM8D+C3gd6MXeJRYCJpH/7tVPIJJnAFSz5P5SVc4I5JOSa0df6KxCYU
U6zzmYS6euac4IhZLXRHUARnbaLtVn6GbbMi1Rx1QbqVaVIHslYFuVIwncyVtbVb
gKrM5RYob7NN1Tz3U+SB9ZQaiT/xI8Go7Tt5hJJGPGXXiHs8R8bUICW67NSlwpmb
w1vXPQmwLxyTuUW6Wj/08Nqjg6t4Oo9pk8/nv39dsg/3aNg1WF4utHgeiKe48s2e
E3q3gvGZDA1MmTDfxFUyfyksEr02V8CYLH+a/5PgW9DIpaPlrhVdB4LX9MZ+8bVj
jtKyqIclmulTUcG0IYWqXD+P7QHWDgO8qyUbKfdTE/OoocTwPD7aZuwnRJWEjz7J
cCYG4IJDGvqG0M0pM7PZ7fwmUZDgXkzLD3JEcaiYLl0kGIUtOuGox8besQb99zv9
dfaHs0/y6cBy4Vmr6FGjVqUyiqr/gnIT76SF2dznotD0J217M8nu4EB1HKnlIXky
9h9xAna/zVsff6w6YyId+yoXDmYa8g48n+II2Eu/NlBtilSJnsHbSC8Am/YiPl6j
XmngalcI3HGRnKr/lC7Gq4b4TguvlMPzpo9I78kl4cZZidZt4WqBAS5jOajASLeW
oELkbrWT9wpUqppaXErCM30m2hHLfhNF2TAXiz+9X5t/t2HicYQocIKmpm/a/wQY
2jw/biTbZpjbEWA/AewQP5rcIaAnU94PsIYqIW3xaT1RLiqxWcThcN+M16I8Na9o
kuoajhqrTh/7RF9W0phdd2+jB67xmqulSOeDAIcf0nvgnEKk65CPy24ZupEjO4to
kjUi655W0EcP8R1RD7pXxOulQwu6RBEXxMuJHjx56lTvxs8SXWqzmk54CiTbWc1l
ksaxVNrUmrioIAk0i2uM0kjPSai2BMbE6XfLGqV+Y3CBJ7pI98mbHNHTkcZA+RsM
8IhZtVBJYsI0bYldPfzfeV1mY6As0eRO4ZuvQtG3IinqWJ2cv3XcXj8jno6O62mI
1x+MJ/I7RLODcXoO/lasg55x7FeR5ht0fHTZClrM0F8LpT75zMobVXDj5Un1TryA
46bVd6t5Z6z6qjusG1YXvUm1VSRGFgo0l95qFS4zqevSzuWDyLeU+CXWg/vM2tg0
yf9q+RB6PClJxoHpk1xpffLJWgzwtEGSJWBHz8I6UqKzipK+a5i4Kwyoaxx2dzUP
VqAVbh1lwNA67OE2tNaBpuvHPOxlV5VjzqJTUtPtIa6xt4zNbhEFvziHLmbG1Ykx
VBuHPI/VacB1eRB0U1W6To58whrX1DHMi02wLjLudEDGAFHseXF/VHgrDzjxpzoC
sk9nALmmhS/KZRUoAyxtpu2pYL7Ztxs5uNFbYv+ooSgjk+HBgxMuDsjyUDBCnH8Z
ZOPeayBbYVJpb5kfyRYH3qkoThJ3OcBTXa1lYubwCY+IM/prk5BFSO6t3aiR7v2h
oJ4ZygydV/MSCCh0hLPr1WNYTf2HqwBcjqxGaPgYjPgGvnTkhJDw596VziCEQoa1
HBNKxDquZprvpHH3O2qNvFtG4YpYpLbA5L4Ex5WhZEM8fzmq5sggDMI80X6H7c/K
4z4sRF0o+TYkvfDLUrbi9GSNG7BBCjp3AltuaFBxbJJfTH08bDf8Vl66ZMYdGMUA
5bjzRXpct2uqL5cdFEzSUThluRQ/iH5nTuNqW6Scp/d2oIiEYTUq+xjBP0hLt4GD
Oskjy/IWOlbVt00v2H/623f+Pc0oGDmTSWSv3nRbFb4Q1snz9kaI3c+n9E4TU5kz
sA7EkE92ixCP8r3W+WBXJGvBeCXZRr17DSYarxw5yUN9sun2Ks6iAUwwc/CnX8qE
SNnJXHcMl08BOm0OUNRyB1X79wyRH8L2at7uwDJ9DsJD3DSg1/T2ZeAH2Ig0T5Va
TPHdv7ibrk23hFVcvpXpGg2BMSRve8LQc7kzR9wkCyhTBwVjvDa5yCP5Ou/jLwga
P2cdQ6m96/DC+lfjUC695ulA7qHcZWdR9dmFfdbjmpaq/rwLrM2qrxX3O0u7CS1X
pykaOSTM9XudK1lGUY+0DgFGZmGyl8U9VwHP8FGirwhx+4bvJy5625zhUWR5kwRq
DsP+E1hug0/lKPkp3wxmgnjL6LJ+MDtIxHXDyW2yiD0BizPYmJp7hYyeguqJ/i6t
TOEsipKzgC6Imosdf9EOio/uEL5ZR+VdT0FU41NdmutEnLydVNfPxNjQBCJnMgyv
mDYsfEInt9LFs+cpN1NVPTgXxWjuU0M67f23GKnqh5ZLzy2dZp6VzMg1FElWw8v6
Faomzs5APL8BXHn76sEaWo+EIXaozjNlJCts+inrVXsh2tVvdmiugzV06Fuqo7+t
a1CIJglf93/MkgwYODtADZl/Sp/XgYkmjONZCuNgTog2DdlVmwW4f4QGNok0u+lk
ZQlX1qyxi8WgKNTcJhE3R1X6UMjSDxDl8U+lSc7/dy9rxzcX8P4p7d0eSn/pr2pb
+/3YFYrhlguRPf3vBCNUsH9TFIzhdBMJ6B/TbnlpprrSfvFwcF5ptPQ9kW/Sg1KC
WtLsA4kyj20XyEGb2OGFKeZ+VRRXg0f0d19c/b9xkCoMaJv805owddD+j1oOnqle
eAPGsnuqzfBy2wyPpdz4vCuqs+lfYTjWN36f2coSBxzbQBGuo+Zt2w97gLudVtig
2C6ti0W1lRHPrk3UsUZS1Z/fuR2tOEGAmJQFk+vXCoDGGRIC7CRV7iRAPJkvBfRj
4PrRE198t5jan00skCx9fgxeBWl27Zh7gIi8PQ1wdQ+7MflQ9WyZXP/VcsfF9PuR
p59WZDIX8NkweGw1Wl8cD6GmLb1tJ59hmVqsUc3owfVGxaPyzeVhXPassKKu582f
VydptXtnlzKEErLhhglqZZanODM6qYlgPRBxc0WWH6ghy43InYlpwwWeZddRXIXo
sa/2x23ssYv15V+MOrtaEpbSJ5yDX3rMo1Rv04aUUrCpE8R+Ho802i+6BBGFnGVn
k/iBMJF1OP4ucZSWHeXRL+EOIzclyJtHXbXhQNl7qz3urlfMOLKvjxSmK2vYZNG/
oZ8FAXvvm/JLbSXMJo7dXgdZ67ixoy3HIRaldj0plHPBya8wc/10a1UJx+URo+Fv
mDxPb9075VveLlkPVBQn8rYAE/Xp1lk17XqPSQN+Wu81kLTyBg0ewBC5DYzOPuaZ
Sj7M93sdaAQK7tT/SKxZ9eYTywfSH8H5xlGSEmIQH9e4EtAQ2tVYXoe826EQ2d6D
RVESZ8GDND/Gl7XEX1PCoPIC8IIUoqv5hul9FM1szxUv56YLXMJNA+fhRVLQevWe
G8qUxpsZgxrHp6KTNlinjgAM7l8F0+3Nhesxg7/j9qOTmpAPgx9YI4To1k1OLcKz
RkbtZ4bxsoQGk6jXosf6vQmPgU2cWFCTgtHyTfbChLaz9VxKf81X6P+w4X2o1fUW
rT0Sa08IKmX74opeFksPEIFrSBHC+37DCzt8Upz8GuR0LV/pm3oJsTdiqHhHw2R8
3wrahx49TSzb52Rn3aB0nlKCzIbRrzlfH+KRkXEgM/xLabTBXgHJOCOB0sFHh6dX
jmuQb6asulXTZRHuZba1s1DNDr4XlntHGZzfZQZJJE/bzVVZqWdq7RD/MsL5hXHA
YDP1GN4lND5CGLLoVhzDRckGoVJ2J3OSDAXDMn+Cmr0=
//pragma protect end_data_block
//pragma protect digest_block
zXKPSnPslyE3OdH5nmd6nMJ6pcs=
//pragma protect end_digest_block
//pragma protect end_protected
