// Copyright (C) 2019  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 19.1.0 Build 670 09/22/2019 SJ Lite Edition"

// DATE "11/26/2019 18:26:51"

// 
// Device: Altera 10M08SAE144C8G Package EQFP144
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module cic (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	in_error,
	in_valid,
	in_ready,
	in0_data,
	in1_data,
	in2_data,
	in3_data,
	in4_data,
	in5_data,
	in6_data,
	in7_data,
	in8_data,
	out_data,
	out_error,
	out_valid,
	out_ready,
	out_startofpacket,
	out_endofpacket,
	out_channel,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	[1:0] in_error;
input 	in_valid;
output 	in_ready;
input 	[0:0] in0_data;
input 	[0:0] in1_data;
input 	[0:0] in2_data;
input 	[0:0] in3_data;
input 	[0:0] in4_data;
input 	[0:0] in5_data;
input 	[0:0] in6_data;
input 	[0:0] in7_data;
input 	[0:0] in8_data;
output 	[18:0] out_data;
output 	[1:0] out_error;
output 	out_valid;
input 	out_ready;
output 	out_startofpacket;
output 	out_endofpacket;
output 	[3:0] out_channel;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \cic_ii_0|core|input_sink|sink_FIFO|auto_generated|dpfifo|full_dff~q ;
wire \cic_ii_0|core|output_source_1|source_valid_s~q ;
wire \cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ;
wire \cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \cic_ii_0|out_data[0]~combout ;
wire \cic_ii_0|out_data[1]~combout ;
wire \cic_ii_0|out_data[2]~combout ;
wire \cic_ii_0|out_data[3]~combout ;
wire \cic_ii_0|out_data[4]~combout ;
wire \cic_ii_0|out_data[5]~combout ;
wire \cic_ii_0|out_data[6]~combout ;
wire \cic_ii_0|out_data[7]~combout ;
wire \cic_ii_0|out_data[8]~combout ;
wire \cic_ii_0|out_data[9]~combout ;
wire \cic_ii_0|out_data[10]~combout ;
wire \cic_ii_0|out_data[11]~combout ;
wire \cic_ii_0|out_data[12]~combout ;
wire \cic_ii_0|out_data[13]~combout ;
wire \cic_ii_0|out_data[14]~combout ;
wire \cic_ii_0|out_data[15]~combout ;
wire \cic_ii_0|out_data[16]~combout ;
wire \cic_ii_0|out_data[17]~combout ;
wire \cic_ii_0|out_data[18]~combout ;
wire \cic_ii_0|core|output_source_1|Equal0~0_combout ;
wire \cic_ii_0|core|output_source_1|Equal1~0_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ;
wire \clk~input_o ;
wire \in_valid~input_o ;
wire \reset_n~input_o ;
wire \out_ready~input_o ;
wire \in5_data[0]~input_o ;
wire \in6_data[0]~input_o ;
wire \in4_data[0]~input_o ;
wire \in7_data[0]~input_o ;
wire \in2_data[0]~input_o ;
wire \in1_data[0]~input_o ;
wire \in0_data[0]~input_o ;
wire \in3_data[0]~input_o ;
wire \in8_data[0]~input_o ;
wire \in_error[0]~input_o ;
wire \in_error[1]~input_o ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TCKUTAP ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|AMGP4450_0~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:1:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:2:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:3:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:4:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:5:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:6:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:7:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:8:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:9:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:10:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:11:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:12:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:13:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_0~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_1~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_1~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_2~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_2~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_3~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_3~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_4~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_4~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_5~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_5~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_6~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_6~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~15_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[10]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~16_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[11]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~17_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[12]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal12~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~18_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[13]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~14_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[14]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~20_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[15]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~2_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~19_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[16]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~13_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[17]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~12_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~3_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~4_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~5_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~6_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~11_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~10_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[2]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~9_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[3]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal3~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~8_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[4]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~7_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[5]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~6_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[6]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal6~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~5_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[7]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~4_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[8]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~3_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[9]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~2_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[18]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ;
wire \~GND~combout ;
wire \altera_internal_jtag~TDIUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal2~1_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~1_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~3_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~4_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~5_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[3]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Equal3~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~8_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[4]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~9_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[5]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Equal5~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~10_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~11_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[7]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~12_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~13_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[8]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Equal8~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~6_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[9]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~7_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[10]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~4_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~2_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[11]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~2_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~3_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ;
wire \nabboc|pzdyqx_impl_inst|BWHK8171_1~q ;
wire \nabboc|pzdyqx_impl_inst|BWHK8171_2~q ;
wire \nabboc|pzdyqx_impl_inst|process_0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ;
wire \nabboc|pzdyqx_impl_inst|process_0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|FWCA1915[3]~q ;
wire \nabboc|pzdyqx_impl_inst|ZIVV0726~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ZIVV0726~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal2~2_combout ;
wire \nabboc|pzdyqx_impl_inst|FWCA1915[2]~q ;
wire \nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ;
wire \nabboc|pzdyqx_impl_inst|NJQG9082~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~23_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~15 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~22_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~10 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~12 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~14 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~6 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~20_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8_combout ;
wire \nabboc|pzdyqx_impl_inst|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal2~0_combout ;
wire \nabboc|pzdyqx_impl_inst|FWCA1915[1]~q ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~3_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~1_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~1 ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~2_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~2_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~3 ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~4_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~q ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~5 ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~6_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~q ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~7 ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~8_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~0_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4]~q ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~4_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[0]~0_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~5_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~6_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[1]~1_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~7_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[2]~2_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~8_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~9_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[3]~3_combout ;
wire \nabboc|pzdyqx_impl_inst|comb~0_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[3]~q ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[2]~q ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[1]~q ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[0]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~12_combout ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[12]~q ;
wire \nabboc|pzdyqx_impl_inst|dr_scan~combout ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~11_combout ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[11]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~10_combout ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[10]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~9_combout ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[9]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~8_combout ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[8]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~7_combout ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[7]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~6_combout ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[6]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~5_combout ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[5]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~4_combout ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[4]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~3_combout ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[3]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~2_combout ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[2]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~1_combout ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[1]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~0_combout ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[0]~q ;
wire \nabboc|pzdyqx_impl_inst|tdo~0_combout ;
wire \nabboc|pzdyqx_impl_inst|KNOR6738~q ;
wire \nabboc|pzdyqx_impl_inst|tdo~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ;
wire \altera_internal_jtag~TDO ;


cic_cic_cic_ii_0 cic_ii_0(
	.full_dff(\cic_ii_0|core|input_sink|sink_FIFO|auto_generated|dpfifo|full_dff~q ),
	.source_valid_s(\cic_ii_0|core|output_source_1|source_valid_s~q ),
	.q_b_22(\cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ),
	.q_b_19(\cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.q_b_20(\cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.q_b_21(\cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.out_data_0(\cic_ii_0|out_data[0]~combout ),
	.out_data_1(\cic_ii_0|out_data[1]~combout ),
	.out_data_2(\cic_ii_0|out_data[2]~combout ),
	.out_data_3(\cic_ii_0|out_data[3]~combout ),
	.out_data_4(\cic_ii_0|out_data[4]~combout ),
	.out_data_5(\cic_ii_0|out_data[5]~combout ),
	.out_data_6(\cic_ii_0|out_data[6]~combout ),
	.out_data_7(\cic_ii_0|out_data[7]~combout ),
	.out_data_8(\cic_ii_0|out_data[8]~combout ),
	.out_data_9(\cic_ii_0|out_data[9]~combout ),
	.out_data_10(\cic_ii_0|out_data[10]~combout ),
	.out_data_11(\cic_ii_0|out_data[11]~combout ),
	.out_data_12(\cic_ii_0|out_data[12]~combout ),
	.out_data_13(\cic_ii_0|out_data[13]~combout ),
	.out_data_14(\cic_ii_0|out_data[14]~combout ),
	.out_data_15(\cic_ii_0|out_data[15]~combout ),
	.out_data_16(\cic_ii_0|out_data[16]~combout ),
	.out_data_17(\cic_ii_0|out_data[17]~combout ),
	.out_data_18(\cic_ii_0|out_data[18]~combout ),
	.Equal0(\cic_ii_0|core|output_source_1|Equal0~0_combout ),
	.Equal1(\cic_ii_0|core|output_source_1|Equal1~0_combout ),
	.GND_port(\~GND~combout ),
	.NJQG9082(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.clk(\clk~input_o ),
	.in_valid(\in_valid~input_o ),
	.reset_n(\reset_n~input_o ),
	.out_ready(\out_ready~input_o ),
	.in5_data_0(\in5_data[0]~input_o ),
	.in6_data_0(\in6_data[0]~input_o ),
	.in4_data_0(\in4_data[0]~input_o ),
	.in7_data_0(\in7_data[0]~input_o ),
	.in2_data_0(\in2_data[0]~input_o ),
	.in1_data_0(\in1_data[0]~input_o ),
	.in0_data_0(\in0_data[0]~input_o ),
	.in3_data_0(\in3_data[0]~input_o ),
	.in8_data_0(\in8_data[0]~input_o ));

assign \clk~input_o  = clk;

assign \in_valid~input_o  = in_valid;

assign \reset_n~input_o  = reset_n;

assign \out_ready~input_o  = out_ready;

assign \in5_data[0]~input_o  = in5_data[0];

assign \in6_data[0]~input_o  = in6_data[0];

assign \in4_data[0]~input_o  = in4_data[0];

assign \in7_data[0]~input_o  = in7_data[0];

assign \in2_data[0]~input_o  = in2_data[0];

assign \in1_data[0]~input_o  = in1_data[0];

assign \in0_data[0]~input_o  = in0_data[0];

assign \in3_data[0]~input_o  = in3_data[0];

assign \in8_data[0]~input_o  = in8_data[0];

assign in_ready = ~ \cic_ii_0|core|input_sink|sink_FIFO|auto_generated|dpfifo|full_dff~q ;

assign out_data[0] = \cic_ii_0|out_data[0]~combout ;

assign out_data[1] = \cic_ii_0|out_data[1]~combout ;

assign out_data[2] = \cic_ii_0|out_data[2]~combout ;

assign out_data[3] = \cic_ii_0|out_data[3]~combout ;

assign out_data[4] = \cic_ii_0|out_data[4]~combout ;

assign out_data[5] = \cic_ii_0|out_data[5]~combout ;

assign out_data[6] = \cic_ii_0|out_data[6]~combout ;

assign out_data[7] = \cic_ii_0|out_data[7]~combout ;

assign out_data[8] = \cic_ii_0|out_data[8]~combout ;

assign out_data[9] = \cic_ii_0|out_data[9]~combout ;

assign out_data[10] = \cic_ii_0|out_data[10]~combout ;

assign out_data[11] = \cic_ii_0|out_data[11]~combout ;

assign out_data[12] = \cic_ii_0|out_data[12]~combout ;

assign out_data[13] = \cic_ii_0|out_data[13]~combout ;

assign out_data[14] = \cic_ii_0|out_data[14]~combout ;

assign out_data[15] = \cic_ii_0|out_data[15]~combout ;

assign out_data[16] = \cic_ii_0|out_data[16]~combout ;

assign out_data[17] = \cic_ii_0|out_data[17]~combout ;

assign out_data[18] = \cic_ii_0|out_data[18]~combout ;

assign out_error[0] = \in_error[0]~input_o ;

assign out_error[1] = \in_error[1]~input_o ;

assign out_valid = \cic_ii_0|core|output_source_1|source_valid_s~q ;

assign out_startofpacket = \cic_ii_0|core|output_source_1|Equal0~0_combout ;

assign out_endofpacket = \cic_ii_0|core|output_source_1|Equal1~0_combout ;

assign out_channel[0] = \cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[19] ;

assign out_channel[1] = \cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[20] ;

assign out_channel[2] = \cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[21] ;

assign out_channel[3] = \cic_ii_0|core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[22] ;

assign altera_reserved_tdo = \altera_internal_jtag~TDO ;

assign \in_error[0]~input_o  = in_error[0];

assign \in_error[1]~input_o  = in_error[1];

assign \altera_reserved_tms~input_o  = altera_reserved_tms;

assign \altera_reserved_tck~input_o  = altera_reserved_tck;

assign \altera_reserved_tdi~input_o  = altera_reserved_tdi;

fiftyfivenm_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdouser(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|AMGP4450_0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:13:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|AMGP4450_0~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|AMGP4450_0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|AMGP4450_0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:1:AMGP4450_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|AMGP4450_0~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:1:AMGP4450_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:1:AMGP4450_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:1:AMGP4450_1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:2:AMGP4450_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:1:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:2:AMGP4450_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:2:AMGP4450_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:2:AMGP4450_1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:3:AMGP4450_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:2:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:3:AMGP4450_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:3:AMGP4450_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:3:AMGP4450_1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:4:AMGP4450_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:3:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:4:AMGP4450_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:4:AMGP4450_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:4:AMGP4450_1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:5:AMGP4450_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:4:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:5:AMGP4450_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:5:AMGP4450_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:5:AMGP4450_1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:6:AMGP4450_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:5:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:6:AMGP4450_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:6:AMGP4450_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:6:AMGP4450_1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:7:AMGP4450_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:6:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:7:AMGP4450_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:7:AMGP4450_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:7:AMGP4450_1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:8:AMGP4450_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:7:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:8:AMGP4450_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:8:AMGP4450_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:8:AMGP4450_1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:9:AMGP4450_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:8:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:9:AMGP4450_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:9:AMGP4450_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:9:AMGP4450_1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:10:AMGP4450_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:9:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:10:AMGP4450_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:10:AMGP4450_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:10:AMGP4450_1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:11:AMGP4450_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:10:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:11:AMGP4450_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:11:AMGP4450_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:11:AMGP4450_1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:12:AMGP4450_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:11:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:12:AMGP4450_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:12:AMGP4450_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:12:AMGP4450_1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:13:AMGP4450_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:12:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:13:AMGP4450_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:13:AMGP4450_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:13:AMGP4450_1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_0~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_0~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_0~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_0~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_0~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_0 (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|SQHZ7915:13:AMGP4450_1~combout ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_0~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_0 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_0 .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_1~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_1~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_1~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_1~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_1~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_1 (
	.clk(!\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_0~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_1~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_1 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_1 .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_2~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_2~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_2~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_2~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_2~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_2 (
	.clk(!\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_1~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_2~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_2 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_2 .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_3~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_3~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_3~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_3~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_3~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_3 (
	.clk(!\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_2~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_3~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_3 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_3 .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_4~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_4~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_4~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_4~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_4~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_4 (
	.clk(!\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_3~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_4~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_4 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_4 .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_5~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_5~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_5~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_5~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_5~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_5 (
	.clk(!\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_4~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_5~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_5 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_5 .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_6~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_6~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_6~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_6~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_6~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_6 (
	.clk(!\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_5~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_6~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_6 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_6 .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7 (
	.clk(!\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_6~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7 .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~15 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[10]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~15_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~15 .lut_mask = 16'h0FF0;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~15 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[10] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[10] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~16 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[11]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[10]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~16_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~16 .lut_mask = 16'hC33C;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~16 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[11] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[11] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~17 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[12]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[10]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[11]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~17_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~17 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~17 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[12] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[12]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[12] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[12] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal12~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[10]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[11]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[12]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal12~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal12~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal12~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~18 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[13]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal12~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~18_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~18 .lut_mask = 16'h0FF0;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~18 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[13] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[13]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[13] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[13] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~14 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[14]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[13]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal12~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~14_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~14 .lut_mask = 16'hC33C;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~14 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[14] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[14]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[14] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[14] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[10]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[11]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[12]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[13]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~20 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[14]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~0_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[15]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~20_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~20 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~20 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[15] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[15]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[15] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[15] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[14]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~2 .lut_mask = 16'hEEEE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~19 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[16]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~2_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[15]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~19_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~19 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~19 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[16] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[16]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[16] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[16] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[14]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~0_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[15]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[16]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~1 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~13 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[17]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~1_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~13_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~13 .lut_mask = 16'hC33C;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~13 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[17] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[17]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[17] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[17] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~12_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~12 .lut_mask = 16'h0FF0;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~12 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~3 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[18]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[2]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~3_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~3 .lut_mask = 16'hFEFF;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~4 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[6]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[5]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~4_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~4 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~5 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[9]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[8]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[7]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~4_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~5_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~5 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~6 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[17]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~1_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~3_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~5_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~6_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~6 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~6 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~11 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~11_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~11 .lut_mask = 16'h7777;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~11 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~10 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[2]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~10_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~10 .lut_mask = 16'hC33C;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~10 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[2] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[2] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~9 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[3]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[2]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~9_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~9 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~9 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[3] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[3] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal3~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[3]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[2]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal3~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal3~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal3~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal3~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~8_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~8 .lut_mask = 16'h0FF0;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~8 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[4] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[4] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~7 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[5]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal3~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~7_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~7 .lut_mask = 16'hC33C;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~7 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[5] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[5] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~6 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[6]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[5]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal3~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~6_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~6 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~6 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[6] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[6] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal6~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[6]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[5]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal3~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal6~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal6~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal6~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[7]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal6~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~5_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~5 .lut_mask = 16'h0FF0;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~5 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[7] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[7] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~4 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[8]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[7]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal6~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~4_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~4 .lut_mask = 16'hC33C;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~4 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[8] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[8] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~3 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[9]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[8]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[7]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal6~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~3_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~3 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~3 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[9] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[9] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[9]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[8]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[7]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal6~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[18]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[17]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~1_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~2 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~2 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[18] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[18]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[18] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[18] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .lut_mask = 16'h0FF0;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .lut_mask = 16'hC33C;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .lut_mask = 16'hFF7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .power_up = "low";

fiftyfivenm_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~GND~combout ),
	.cout());
defparam \~GND .lut_mask = 16'h0000;
defparam \~GND .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .lut_mask = 16'h7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~6 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~10 (
	.dataa(\~GND~combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~6_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~10 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~5 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~10_combout ),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~11 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~11_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~1 .lut_mask = 16'hEEEE;
defparam \nabboc|pzdyqx_impl_inst|Equal2~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~0 .lut_mask = 16'h7777;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~1 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~1 .lut_mask = 16'h3CFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~1 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~3 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~3_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~3 .lut_mask = 16'h96FF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~3 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~4 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[3]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~4_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~4 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~5 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~5_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~5 .lut_mask = 16'hAAFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~5 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[3] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[3] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Equal3~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal3~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal3~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal3~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~8 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[4]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal3~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~8_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~8 .lut_mask = 16'h3CFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~8 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[4] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[4] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~9 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[5]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[4]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal3~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~9_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~9 .lut_mask = 16'h96FF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~9 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[5] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[5] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Equal5~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[4]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[5]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal3~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal5~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal5~0 .lut_mask = 16'hFEFE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal5~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~10 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal5~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~10_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~10 .lut_mask = 16'h3CFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~10 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~11 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[7]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal5~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~11_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~11 .lut_mask = 16'h96FF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~11 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[7] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[7] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~12 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[8]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[7]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal5~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~12_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~12 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~13 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~12_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~13_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~13 .lut_mask = 16'hAAFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~13 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[8] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[8] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Equal8~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[7]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[8]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal5~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal8~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal8~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal8~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~6 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[9]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal8~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~6_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~6 .lut_mask = 16'h3CFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~6 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[9] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[9] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~7 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[10]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[9]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal8~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~7_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~7 .lut_mask = 16'h96FF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~7 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[10] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[10] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~4 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[9]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~4_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~4 .lut_mask = 16'hEEEE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[11]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~4_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal8~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~2 .lut_mask = 16'h96FF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~2 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[11] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[11] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[11]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~1 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[9]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[10]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[4]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~1 .lut_mask = 16'hEFFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[5]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[7]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[8]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~2 .lut_mask = 16'h7FFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~3 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~1_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~3_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~3 .lut_mask = 16'hFEFE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~3 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|BWHK8171_1 (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|BWHK8171_1~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|BWHK8171_1 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|BWHK8171_1 .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|BWHK8171_2 (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|BWHK8171_1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|BWHK8171_2~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|BWHK8171_2 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|BWHK8171_2 .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|process_0~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|FWCA1915[3]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|BWHK8171_2~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|process_0~0 .lut_mask = 16'hEEEE;
defparam \nabboc|pzdyqx_impl_inst|process_0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .lut_mask = 16'hEFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 .lut_mask = 16'hFDFD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~6 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~6_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~7 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~5_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~6_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~12 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~12_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13 .lut_mask = 16'hACFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~7 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~7_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~14 .lut_mask = 16'hFFAC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~14 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~14_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3 .lut_mask = 16'hEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .lut_mask = 16'hB8FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|process_0~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|FWCA1915[2]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|process_0~1 .lut_mask = 16'hFEFF;
defparam \nabboc|pzdyqx_impl_inst|process_0~1 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|FWCA1915[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~1_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|FWCA1915[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|FWCA1915[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|FWCA1915[3] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|ZIVV0726~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|ZIVV0726~q ),
	.datab(\nabboc|pzdyqx_impl_inst|FWCA1915[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ZIVV0726~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ZIVV0726~0 .lut_mask = 16'hEEEE;
defparam \nabboc|pzdyqx_impl_inst|ZIVV0726~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ZIVV0726 (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ZIVV0726~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|BWHK8171_2~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ZIVV0726~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ZIVV0726 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ZIVV0726 .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8 (
	.dataa(\nabboc|pzdyqx_impl_inst|ZIVV0726~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~14_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~0 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4 .lut_mask = 16'h0FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~2 .lut_mask = 16'hAAFF;
defparam \nabboc|pzdyqx_impl_inst|Equal2~2 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|FWCA1915[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~2_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|FWCA1915[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|FWCA1915[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|FWCA1915[2] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|NJQG9082~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.datab(\nabboc|pzdyqx_impl_inst|FWCA1915[2]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|BWHK8171_1~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ZIVV0726~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|NJQG9082~0 .lut_mask = 16'hFEFF;
defparam \nabboc|pzdyqx_impl_inst|NJQG9082~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|NJQG9082 (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_ZNXJ5711_gen_0:cycloneiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|NJQG9082 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|NJQG9082 .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 (
	.dataa(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~14_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 .lut_mask = 16'h55AA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~15 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~23 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~23_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~23 .lut_mask = 16'hFFFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~23 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~15 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 .lut_mask = 16'h5AAF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 .lut_mask = 16'h5A5A;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~13 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~22 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~13_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~22_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~22 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~22 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 .lut_mask = 16'h6FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .lut_mask = 16'hD8FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~6 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5 .lut_mask = 16'h55AA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~6 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~9_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~10 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~9 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~9 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~10 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~12 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11 .lut_mask = 16'h5AAF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~8 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~8 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~7_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~8_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~12 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~14 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~7_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~8_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~14 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15 .lut_mask = 16'h5A5A;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~7_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~8_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~7 .lut_mask = 16'hFFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~7_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~8_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~7_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~8_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~20 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~20_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~20 .lut_mask = 16'hDFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~20 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~8 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~8_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~9 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~20_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 .lut_mask = 16'hEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 .lut_mask = 16'h0C3F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17 .lut_mask = 16'hEDDE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18 .lut_mask = 16'hD77D;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15 .lut_mask = 16'hEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16 .lut_mask = 16'hDF8F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .lut_mask = 16'h0FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena .lut_mask = 16'hFFFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|Equal0~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal0~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|Equal0~0 .lut_mask = 16'h7777;
defparam \nabboc|pzdyqx_impl_inst|Equal0~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|FWCA1915[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal0~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|FWCA1915[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|FWCA1915[0] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~0 .lut_mask = 16'hAAFF;
defparam \nabboc|pzdyqx_impl_inst|Equal2~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|FWCA1915[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|FWCA1915[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|FWCA1915[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|FWCA1915[1] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|Add0~0_combout ),
	.cout(\nabboc|pzdyqx_impl_inst|VWQM3427|Add0~1 ));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~0 .lut_mask = 16'h55AA;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|Equal0~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|Equal0~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|Equal0~0 .lut_mask = 16'hEFFF;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|Equal0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~3 (
	.dataa(\nabboc|pzdyqx_impl_inst|VWQM3427|Add0~0_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|VWQM3427|Equal0~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~3_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~3 .lut_mask = 16'h9966;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0 .lut_mask = 16'hEEEE;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~1 .lut_mask = 16'hEFFF;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~1 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~3_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nabboc|pzdyqx_impl_inst|VWQM3427|Add0~1 ),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|Add0~2_combout ),
	.cout(\nabboc|pzdyqx_impl_inst|VWQM3427|Add0~3 ));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~2 .lut_mask = 16'h5A5F;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|VWQM3427|Add0~2_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|VWQM3427|Equal0~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~2 .lut_mask = 16'h9966;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~2 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~2_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~4 (
	.dataa(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nabboc|pzdyqx_impl_inst|VWQM3427|Add0~3 ),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|Add0~4_combout ),
	.cout(\nabboc|pzdyqx_impl_inst|VWQM3427|Add0~5 ));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~4 .lut_mask = 16'h5AAF;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~4 .sum_lutc_input = "cin";

dffeas \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|VWQM3427|Add0~4_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~6 (
	.dataa(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nabboc|pzdyqx_impl_inst|VWQM3427|Add0~5 ),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|Add0~6_combout ),
	.cout(\nabboc|pzdyqx_impl_inst|VWQM3427|Add0~7 ));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~6 .lut_mask = 16'h5A5F;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~6 .sum_lutc_input = "cin";

dffeas \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|VWQM3427|Add0~6_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~8 (
	.dataa(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\nabboc|pzdyqx_impl_inst|VWQM3427|Add0~7 ),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|Add0~8_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~8 .lut_mask = 16'h5A5A;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|Add0~8 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|VWQM3427|Add0~8_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|VWQM3427|Equal0~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~0 .lut_mask = 16'h9966;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~4 (
	.dataa(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~4_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~4 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[0]~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~4_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[0]~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[0]~0 .lut_mask = 16'hCC55;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~5 (
	.dataa(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~5_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~5 .lut_mask = 16'hF6F6;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~6 (
	.dataa(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~q ),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~6_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~6 .lut_mask = 16'h66FF;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[1]~1 (
	.dataa(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~5_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~6_combout ),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[1]~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[1]~1 .lut_mask = 16'hAACC;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[1]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~7 (
	.dataa(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~7_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~7 .lut_mask = 16'hEFFF;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[2]~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~7_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~6_combout ),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[2]~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[2]~2 .lut_mask = 16'hAACC;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[2]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~8 (
	.dataa(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~8_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~8 .lut_mask = 16'hF6FF;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~9 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~9_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~9 .lut_mask = 16'hC33C;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[3]~3 (
	.dataa(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~8_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~9_combout ),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[3]~3_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[3]~3 .lut_mask = 16'hAA33;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|comb~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|comb~0 .lut_mask = 16'hFEFF;
defparam \nabboc|pzdyqx_impl_inst|comb~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[3]~3_combout ),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(!\nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[3] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[2]~2_combout ),
	.asdata(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[3]~q ),
	.clrn(!\nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[2] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[1]~1_combout ),
	.asdata(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[2]~q ),
	.clrn(!\nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[1] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[0]~0_combout ),
	.asdata(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[1]~q ),
	.clrn(!\nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[0] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~12_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~12 .lut_mask = 16'hFEFF;
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~12 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[12]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[12] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[12] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|dr_scan (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|dr_scan .lut_mask = 16'hAAFF;
defparam \nabboc|pzdyqx_impl_inst|dr_scan .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~11 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[11]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[12]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~11_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~11 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~11 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[11] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~10 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[10]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[11]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~10_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~10 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~10 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[10] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~9 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[9]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[10]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~9_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~9 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~9 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[9] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~8 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[8]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[9]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~8_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~8 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~8 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[8] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~7 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[7]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~7_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~7 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~7 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[7] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~6 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[7]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~6_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~6 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~6 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[6] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~5 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[5]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[6]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~5_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~5 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~5 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[5] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~4 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[4]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~4_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~4 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~4 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[4] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~3 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[3]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~3_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~3 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~3 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[3] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~2 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~2 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[2] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~1 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~1 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~1 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[1] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~0 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[0] .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|tdo~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|FWCA1915[1]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|tdo~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|tdo~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|tdo~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|KNOR6738 (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|KNOR6738~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|KNOR6738 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|KNOR6738 .power_up = "low";

fiftyfivenm_lcell_comb \nabboc|pzdyqx_impl_inst|tdo~1 (
	.dataa(\nabboc|pzdyqx_impl_inst|tdo~0_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|KNOR6738~q ),
	.datac(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|FWCA1915[1]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|tdo~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|tdo~1 .lut_mask = 16'hEFFF;
defparam \nabboc|pzdyqx_impl_inst|tdo~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|tdo~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo (
	.clk(!\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|~GND~combout ),
	.cout());
defparam \auto_hub|~GND .lut_mask = 16'h0000;
defparam \auto_hub|~GND .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .sum_lutc_input = "datac";

endmodule

module cic_cic_cic_ii_0 (
	full_dff,
	source_valid_s,
	q_b_22,
	q_b_19,
	q_b_20,
	q_b_21,
	out_data_0,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_5,
	out_data_6,
	out_data_7,
	out_data_8,
	out_data_9,
	out_data_10,
	out_data_11,
	out_data_12,
	out_data_13,
	out_data_14,
	out_data_15,
	out_data_16,
	out_data_17,
	out_data_18,
	Equal0,
	Equal1,
	GND_port,
	NJQG9082,
	clk,
	in_valid,
	reset_n,
	out_ready,
	in5_data_0,
	in6_data_0,
	in4_data_0,
	in7_data_0,
	in2_data_0,
	in1_data_0,
	in0_data_0,
	in3_data_0,
	in8_data_0)/* synthesis synthesis_greybox=1 */;
output 	full_dff;
output 	source_valid_s;
output 	q_b_22;
output 	q_b_19;
output 	q_b_20;
output 	q_b_21;
output 	out_data_0;
output 	out_data_1;
output 	out_data_2;
output 	out_data_3;
output 	out_data_4;
output 	out_data_5;
output 	out_data_6;
output 	out_data_7;
output 	out_data_8;
output 	out_data_9;
output 	out_data_10;
output 	out_data_11;
output 	out_data_12;
output 	out_data_13;
output 	out_data_14;
output 	out_data_15;
output 	out_data_16;
output 	out_data_17;
output 	out_data_18;
output 	Equal0;
output 	Equal1;
input 	GND_port;
input 	NJQG9082;
input 	clk;
input 	in_valid;
input 	reset_n;
input 	out_ready;
input 	in5_data_0;
input 	in6_data_0;
input 	in4_data_0;
input 	in7_data_0;
input 	in2_data_0;
input 	in1_data_0;
input 	in0_data_0;
input 	in3_data_0;
input 	in8_data_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;


cic_alt_cic_core core(
	.full_dff(full_dff),
	.q_b_0(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_1(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_2(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_4(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_5(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_6(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_7(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_8(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.q_b_9(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.q_b_10(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.q_b_11(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.q_b_12(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.q_b_13(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.q_b_14(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.q_b_15(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.q_b_16(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.q_b_17(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.q_b_18(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.source_valid_s(source_valid_s),
	.q_b_22(q_b_22),
	.q_b_19(q_b_19),
	.q_b_20(q_b_20),
	.q_b_21(q_b_21),
	.Equal0(Equal0),
	.Equal1(Equal1),
	.GND_port(GND_port),
	.clk(clk),
	.in_valid(in_valid),
	.reset_n(reset_n),
	.out_ready(out_ready),
	.in5_data_0(in5_data_0),
	.in6_data_0(in6_data_0),
	.in4_data_0(in4_data_0),
	.in7_data_0(in7_data_0),
	.in2_data_0(in2_data_0),
	.in1_data_0(in1_data_0),
	.in0_data_0(in0_data_0),
	.in3_data_0(in3_data_0),
	.in8_data_0(in8_data_0));

fiftyfivenm_lcell_comb \out_data[0] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_0),
	.cout());
defparam \out_data[0] .lut_mask = 16'hAAFF;
defparam \out_data[0] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[1] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_1),
	.cout());
defparam \out_data[1] .lut_mask = 16'hAAFF;
defparam \out_data[1] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[2] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_2),
	.cout());
defparam \out_data[2] .lut_mask = 16'hAAFF;
defparam \out_data[2] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[3] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_3),
	.cout());
defparam \out_data[3] .lut_mask = 16'hAAFF;
defparam \out_data[3] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[4] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_4),
	.cout());
defparam \out_data[4] .lut_mask = 16'hAAFF;
defparam \out_data[4] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[5] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_5),
	.cout());
defparam \out_data[5] .lut_mask = 16'hAAFF;
defparam \out_data[5] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[6] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_6),
	.cout());
defparam \out_data[6] .lut_mask = 16'hAAFF;
defparam \out_data[6] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[7] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_7),
	.cout());
defparam \out_data[7] .lut_mask = 16'hAAFF;
defparam \out_data[7] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[8] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_8),
	.cout());
defparam \out_data[8] .lut_mask = 16'hAAFF;
defparam \out_data[8] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[9] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_9),
	.cout());
defparam \out_data[9] .lut_mask = 16'hAAFF;
defparam \out_data[9] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[10] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_10),
	.cout());
defparam \out_data[10] .lut_mask = 16'hAAFF;
defparam \out_data[10] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[11] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_11),
	.cout());
defparam \out_data[11] .lut_mask = 16'hAAFF;
defparam \out_data[11] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[12] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_12),
	.cout());
defparam \out_data[12] .lut_mask = 16'hAAFF;
defparam \out_data[12] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[13] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_13),
	.cout());
defparam \out_data[13] .lut_mask = 16'hAAFF;
defparam \out_data[13] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[14] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_14),
	.cout());
defparam \out_data[14] .lut_mask = 16'hAAFF;
defparam \out_data[14] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[15] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_15),
	.cout());
defparam \out_data[15] .lut_mask = 16'hAAFF;
defparam \out_data[15] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[16] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_16),
	.cout());
defparam \out_data[16] .lut_mask = 16'hAAFF;
defparam \out_data[16] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[17] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_17),
	.cout());
defparam \out_data[17] .lut_mask = 16'hAAFF;
defparam \out_data[17] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[18] (
	.dataa(\core|output_source_1|source_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(out_data_18),
	.cout());
defparam \out_data[18] .lut_mask = 16'hAAFF;
defparam \out_data[18] .sum_lutc_input = "datac";

endmodule

module cic_alt_cic_core (
	full_dff,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	source_valid_s,
	q_b_22,
	q_b_19,
	q_b_20,
	q_b_21,
	Equal0,
	Equal1,
	GND_port,
	clk,
	in_valid,
	reset_n,
	out_ready,
	in5_data_0,
	in6_data_0,
	in4_data_0,
	in7_data_0,
	in2_data_0,
	in1_data_0,
	in0_data_0,
	in3_data_0,
	in8_data_0)/* synthesis synthesis_greybox=1 */;
output 	full_dff;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	source_valid_s;
output 	q_b_22;
output 	q_b_19;
output 	q_b_20;
output 	q_b_21;
output 	Equal0;
output 	Equal1;
input 	GND_port;
input 	clk;
input 	in_valid;
input 	reset_n;
input 	out_ready;
input 	in5_data_0;
input 	in6_data_0;
input 	in4_data_0;
input 	in7_data_0;
input 	in2_data_0;
input 	in1_data_0;
input 	in0_data_0;
input 	in3_data_0;
input 	in8_data_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \input_sink|sink_FIFO|auto_generated|dffe_nae~q ;
wire \output_source_1|source_FIFO|auto_generated|dffe_af~q ;
wire \dec_mul|state[0]~q ;
wire \dec_mul|stage_diff[2].auk_dsp_diff|dout[0]~q ;
wire \dec_mul|stage_diff[2].auk_dsp_diff|dout[1]~q ;
wire \dec_mul|stage_diff[2].auk_dsp_diff|dout[2]~q ;
wire \dec_mul|stage_diff[2].auk_dsp_diff|dout[3]~q ;
wire \dec_mul|stage_diff[2].auk_dsp_diff|dout[4]~q ;
wire \dec_mul|stage_diff[2].auk_dsp_diff|dout[5]~q ;
wire \dec_mul|stage_diff[2].auk_dsp_diff|dout[6]~q ;
wire \dec_mul|stage_diff[2].auk_dsp_diff|dout[7]~q ;
wire \dec_mul|stage_diff[2].auk_dsp_diff|dout[8]~q ;
wire \dec_mul|stage_diff[2].auk_dsp_diff|dout[9]~q ;
wire \dec_mul|stage_diff[2].auk_dsp_diff|dout[10]~q ;
wire \dec_mul|stage_diff[2].auk_dsp_diff|dout[11]~q ;
wire \dec_mul|stage_diff[2].auk_dsp_diff|dout[12]~q ;
wire \dec_mul|stage_diff[2].auk_dsp_diff|dout[13]~q ;
wire \dec_mul|stage_diff[2].auk_dsp_diff|dout[14]~q ;
wire \dec_mul|stage_diff[2].auk_dsp_diff|dout[15]~q ;
wire \dec_mul|stage_diff[2].auk_dsp_diff|dout[16]~q ;
wire \dec_mul|stage_diff[2].auk_dsp_diff|dout[17]~q ;
wire \dec_mul|stage_diff[2].auk_dsp_diff|dout[18]~q ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \avalon_controller|ready_FIFO|usedw_process~2_combout ;
wire \avalon_controller|sink_ready_ctrl~1_combout ;
wire \avalon_controller|sink_ready_ctrl~2_combout ;
wire \avalon_controller|stall_reg~q ;
wire \dec_mul|stage_diff[2].auk_dsp_diff|dout_valid~q ;
wire \dec_mul|channel_out_int[3]~q ;
wire \dec_mul|channel_out_int[0]~q ;
wire \dec_mul|channel_out_int[1]~q ;
wire \dec_mul|channel_out_int[2]~q ;


cic_auk_dspip_avalon_streaming_sink input_sink(
	.full_dff(full_dff),
	.dffe_nae(\input_sink|sink_FIFO|auto_generated|dffe_nae~q ),
	.dffe_af(\output_source_1|source_FIFO|auto_generated|dffe_af~q ),
	.data({\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ,\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ,
\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] }),
	.usedw_process(\avalon_controller|ready_FIFO|usedw_process~2_combout ),
	.sink_ready_ctrl(\avalon_controller|sink_ready_ctrl~1_combout ),
	.sink_ready_ctrl1(\avalon_controller|sink_ready_ctrl~2_combout ),
	.GND_port(GND_port),
	.clk(clk),
	.in_valid(in_valid),
	.reset_n(reset_n),
	.at_sink_data({in8_data_0,in7_data_0,in6_data_0,in5_data_0,in4_data_0,in3_data_0,in2_data_0,in1_data_0,in0_data_0}));

cic_alt_cic_dec_miso dec_mul(
	.state_0(\dec_mul|state[0]~q ),
	.dout_0(\dec_mul|stage_diff[2].auk_dsp_diff|dout[0]~q ),
	.dout_1(\dec_mul|stage_diff[2].auk_dsp_diff|dout[1]~q ),
	.dout_2(\dec_mul|stage_diff[2].auk_dsp_diff|dout[2]~q ),
	.dout_3(\dec_mul|stage_diff[2].auk_dsp_diff|dout[3]~q ),
	.dout_4(\dec_mul|stage_diff[2].auk_dsp_diff|dout[4]~q ),
	.dout_5(\dec_mul|stage_diff[2].auk_dsp_diff|dout[5]~q ),
	.dout_6(\dec_mul|stage_diff[2].auk_dsp_diff|dout[6]~q ),
	.dout_7(\dec_mul|stage_diff[2].auk_dsp_diff|dout[7]~q ),
	.dout_8(\dec_mul|stage_diff[2].auk_dsp_diff|dout[8]~q ),
	.dout_9(\dec_mul|stage_diff[2].auk_dsp_diff|dout[9]~q ),
	.dout_10(\dec_mul|stage_diff[2].auk_dsp_diff|dout[10]~q ),
	.dout_11(\dec_mul|stage_diff[2].auk_dsp_diff|dout[11]~q ),
	.dout_12(\dec_mul|stage_diff[2].auk_dsp_diff|dout[12]~q ),
	.dout_13(\dec_mul|stage_diff[2].auk_dsp_diff|dout[13]~q ),
	.dout_14(\dec_mul|stage_diff[2].auk_dsp_diff|dout[14]~q ),
	.dout_15(\dec_mul|stage_diff[2].auk_dsp_diff|dout[15]~q ),
	.dout_16(\dec_mul|stage_diff[2].auk_dsp_diff|dout[16]~q ),
	.dout_17(\dec_mul|stage_diff[2].auk_dsp_diff|dout[17]~q ),
	.dout_18(\dec_mul|stage_diff[2].auk_dsp_diff|dout[18]~q ),
	.q_b_5(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_6(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_4(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_7(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_2(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_1(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_0(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_3(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_8(\input_sink|sink_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.stall_reg(\avalon_controller|stall_reg~q ),
	.dout_valid(\dec_mul|stage_diff[2].auk_dsp_diff|dout_valid~q ),
	.channel_out_int_3(\dec_mul|channel_out_int[3]~q ),
	.channel_out_int_0(\dec_mul|channel_out_int[0]~q ),
	.channel_out_int_1(\dec_mul|channel_out_int[1]~q ),
	.channel_out_int_2(\dec_mul|channel_out_int[2]~q ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_avalon_streaming_controller avalon_controller(
	.dffe_nae(\input_sink|sink_FIFO|auto_generated|dffe_nae~q ),
	.dffe_af(\output_source_1|source_FIFO|auto_generated|dffe_af~q ),
	.usedw_process(\avalon_controller|ready_FIFO|usedw_process~2_combout ),
	.sink_ready_ctrl(\avalon_controller|sink_ready_ctrl~1_combout ),
	.sink_ready_ctrl1(\avalon_controller|sink_ready_ctrl~2_combout ),
	.stall_reg1(\avalon_controller|stall_reg~q ),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_avalon_streaming_source output_source_1(
	.at_source_data({q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.source_valid_s1(source_valid_s),
	.at_source_channel({q_b_22,q_b_21,q_b_20,q_b_19}),
	.dffe_af(\output_source_1|source_FIFO|auto_generated|dffe_af~q ),
	.state_0(\dec_mul|state[0]~q ),
	.data({\dec_mul|stage_diff[2].auk_dsp_diff|dout[18]~q ,\dec_mul|stage_diff[2].auk_dsp_diff|dout[17]~q ,\dec_mul|stage_diff[2].auk_dsp_diff|dout[16]~q ,\dec_mul|stage_diff[2].auk_dsp_diff|dout[15]~q ,\dec_mul|stage_diff[2].auk_dsp_diff|dout[14]~q ,
\dec_mul|stage_diff[2].auk_dsp_diff|dout[13]~q ,\dec_mul|stage_diff[2].auk_dsp_diff|dout[12]~q ,\dec_mul|stage_diff[2].auk_dsp_diff|dout[11]~q ,\dec_mul|stage_diff[2].auk_dsp_diff|dout[10]~q ,\dec_mul|stage_diff[2].auk_dsp_diff|dout[9]~q ,
\dec_mul|stage_diff[2].auk_dsp_diff|dout[8]~q ,\dec_mul|stage_diff[2].auk_dsp_diff|dout[7]~q ,\dec_mul|stage_diff[2].auk_dsp_diff|dout[6]~q ,\dec_mul|stage_diff[2].auk_dsp_diff|dout[5]~q ,\dec_mul|stage_diff[2].auk_dsp_diff|dout[4]~q ,
\dec_mul|stage_diff[2].auk_dsp_diff|dout[3]~q ,\dec_mul|stage_diff[2].auk_dsp_diff|dout[2]~q ,\dec_mul|stage_diff[2].auk_dsp_diff|dout[1]~q ,\dec_mul|stage_diff[2].auk_dsp_diff|dout[0]~q }),
	.Equal0(Equal0),
	.Equal1(Equal1),
	.stall_reg(\avalon_controller|stall_reg~q ),
	.dout_valid(\dec_mul|stage_diff[2].auk_dsp_diff|dout_valid~q ),
	.data_count({\dec_mul|channel_out_int[3]~q ,\dec_mul|channel_out_int[2]~q ,\dec_mul|channel_out_int[1]~q ,\dec_mul|channel_out_int[0]~q }),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n),
	.out_ready(out_ready));

endmodule

module cic_alt_cic_dec_miso (
	state_0,
	dout_0,
	dout_1,
	dout_2,
	dout_3,
	dout_4,
	dout_5,
	dout_6,
	dout_7,
	dout_8,
	dout_9,
	dout_10,
	dout_11,
	dout_12,
	dout_13,
	dout_14,
	dout_15,
	dout_16,
	dout_17,
	dout_18,
	q_b_5,
	q_b_6,
	q_b_4,
	q_b_7,
	q_b_2,
	q_b_1,
	q_b_0,
	q_b_3,
	q_b_8,
	stall_reg,
	dout_valid,
	channel_out_int_3,
	channel_out_int_0,
	channel_out_int_1,
	channel_out_int_2,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	state_0;
output 	dout_0;
output 	dout_1;
output 	dout_2;
output 	dout_3;
output 	dout_4;
output 	dout_5;
output 	dout_6;
output 	dout_7;
output 	dout_8;
output 	dout_9;
output 	dout_10;
output 	dout_11;
output 	dout_12;
output 	dout_13;
output 	dout_14;
output 	dout_15;
output 	dout_16;
output 	dout_17;
output 	dout_18;
input 	q_b_5;
input 	q_b_6;
input 	q_b_4;
input 	q_b_7;
input 	q_b_2;
input 	q_b_1;
input 	q_b_0;
input 	q_b_3;
input 	q_b_8;
input 	stall_reg;
output 	dout_valid;
output 	channel_out_int_3;
output 	channel_out_int_0;
output 	channel_out_int_1;
output 	channel_out_int_2;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \stage_diff[1].auk_dsp_diff|dout[0]~q ;
wire \stage_diff[1].auk_dsp_diff|dout[1]~q ;
wire \stage_diff[1].auk_dsp_diff|dout[2]~q ;
wire \stage_diff[1].auk_dsp_diff|dout[3]~q ;
wire \stage_diff[1].auk_dsp_diff|dout[4]~q ;
wire \stage_diff[1].auk_dsp_diff|dout[5]~q ;
wire \stage_diff[1].auk_dsp_diff|dout[6]~q ;
wire \stage_diff[1].auk_dsp_diff|dout[7]~q ;
wire \stage_diff[1].auk_dsp_diff|dout[8]~q ;
wire \stage_diff[1].auk_dsp_diff|dout[9]~q ;
wire \stage_diff[1].auk_dsp_diff|dout[10]~q ;
wire \stage_diff[1].auk_dsp_diff|dout[11]~q ;
wire \stage_diff[1].auk_dsp_diff|dout[12]~q ;
wire \stage_diff[1].auk_dsp_diff|dout[13]~q ;
wire \stage_diff[1].auk_dsp_diff|dout[14]~q ;
wire \stage_diff[1].auk_dsp_diff|dout[15]~q ;
wire \stage_diff[1].auk_dsp_diff|dout[16]~q ;
wire \stage_diff[1].auk_dsp_diff|dout[17]~q ;
wire \stage_diff[1].auk_dsp_diff|dout[18]~q ;
wire \stage_diff[0].auk_dsp_diff|dout[0]~q ;
wire \stage_diff[0].auk_dsp_diff|dout[1]~q ;
wire \stage_diff[0].auk_dsp_diff|dout[2]~q ;
wire \stage_diff[0].auk_dsp_diff|dout[3]~q ;
wire \stage_diff[0].auk_dsp_diff|dout[4]~q ;
wire \stage_diff[0].auk_dsp_diff|dout[5]~q ;
wire \stage_diff[0].auk_dsp_diff|dout[6]~q ;
wire \stage_diff[0].auk_dsp_diff|dout[7]~q ;
wire \stage_diff[0].auk_dsp_diff|dout[8]~q ;
wire \stage_diff[0].auk_dsp_diff|dout[9]~q ;
wire \stage_diff[0].auk_dsp_diff|dout[10]~q ;
wire \stage_diff[0].auk_dsp_diff|dout[11]~q ;
wire \stage_diff[0].auk_dsp_diff|dout[12]~q ;
wire \stage_diff[0].auk_dsp_diff|dout[13]~q ;
wire \stage_diff[0].auk_dsp_diff|dout[14]~q ;
wire \stage_diff[0].auk_dsp_diff|dout[15]~q ;
wire \stage_diff[0].auk_dsp_diff|dout[16]~q ;
wire \stage_diff[0].auk_dsp_diff|dout[17]~q ;
wire \stage_diff[0].auk_dsp_diff|dout[18]~q ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \Mod2|auto_generated|divider|divider|op_24~1 ;
wire \Mod2|auto_generated|divider|divider|op_24~0_combout ;
wire \Mod2|auto_generated|divider|divider|op_23~1 ;
wire \Mod2|auto_generated|divider|divider|op_23~0_combout ;
wire \Mod2|auto_generated|divider|divider|op_23~3 ;
wire \Mod2|auto_generated|divider|divider|op_23~2_combout ;
wire \Mod2|auto_generated|divider|divider|op_23~5 ;
wire \Mod2|auto_generated|divider|divider|op_23~4_combout ;
wire \Mod2|auto_generated|divider|divider|op_23~7 ;
wire \Mod2|auto_generated|divider|divider|op_23~6_combout ;
wire \Mod2|auto_generated|divider|divider|op_23~9_cout ;
wire \Mod2|auto_generated|divider|divider|op_23~10_combout ;
wire \Mod2|auto_generated|divider|divider|op_24~3 ;
wire \Mod2|auto_generated|divider|divider|op_24~2_combout ;
wire \Mod2|auto_generated|divider|divider|op_24~5 ;
wire \Mod2|auto_generated|divider|divider|op_24~4_combout ;
wire \Mod2|auto_generated|divider|divider|op_24~7 ;
wire \Mod2|auto_generated|divider|divider|op_24~6_combout ;
wire \Mod2|auto_generated|divider|divider|op_24~9_cout ;
wire \Mod2|auto_generated|divider|divider|op_24~10_combout ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \ena_sample~q ;
wire \sample_state[0]~q ;
wire \integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[6]~q ;
wire \integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[1]~q ;
wire \integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[2]~q ;
wire \integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[3]~q ;
wire \integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[4]~q ;
wire \integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[0]~q ;
wire \integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[5]~q ;
wire \integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \Mod0|auto_generated|divider|divider|op_5~1 ;
wire \Mod0|auto_generated|divider|divider|op_5~0_combout ;
wire \Mod0|auto_generated|divider|divider|op_1~1 ;
wire \Mod0|auto_generated|divider|divider|op_1~0_combout ;
wire \Mod0|auto_generated|divider|divider|op_1~3 ;
wire \Mod0|auto_generated|divider|divider|op_1~2_combout ;
wire \Mod0|auto_generated|divider|divider|op_1~5 ;
wire \Mod0|auto_generated|divider|divider|op_1~4_combout ;
wire \Mod0|auto_generated|divider|divider|op_1~6_combout ;
wire \Mod0|auto_generated|divider|divider|op_2~1 ;
wire \Mod0|auto_generated|divider|divider|op_2~0_combout ;
wire \Mod0|auto_generated|divider|divider|op_2~3 ;
wire \Mod0|auto_generated|divider|divider|op_2~2_combout ;
wire \Mod0|auto_generated|divider|divider|op_2~5 ;
wire \Mod0|auto_generated|divider|divider|op_2~4_combout ;
wire \Mod0|auto_generated|divider|divider|op_2~7_cout ;
wire \Mod0|auto_generated|divider|divider|op_2~8_combout ;
wire \Mod0|auto_generated|divider|divider|op_3~1 ;
wire \Mod0|auto_generated|divider|divider|op_3~0_combout ;
wire \Mod0|auto_generated|divider|divider|op_3~3 ;
wire \Mod0|auto_generated|divider|divider|op_3~2_combout ;
wire \Mod0|auto_generated|divider|divider|op_3~5 ;
wire \Mod0|auto_generated|divider|divider|op_3~4_combout ;
wire \Mod0|auto_generated|divider|divider|op_3~7_cout ;
wire \Mod0|auto_generated|divider|divider|op_3~8_combout ;
wire \Mod0|auto_generated|divider|divider|op_4~1 ;
wire \Mod0|auto_generated|divider|divider|op_4~0_combout ;
wire \Mod0|auto_generated|divider|divider|op_4~3 ;
wire \Mod0|auto_generated|divider|divider|op_4~2_combout ;
wire \Mod0|auto_generated|divider|divider|op_4~5 ;
wire \Mod0|auto_generated|divider|divider|op_4~4_combout ;
wire \Mod0|auto_generated|divider|divider|op_4~7_cout ;
wire \Mod0|auto_generated|divider|divider|op_4~8_combout ;
wire \Mod0|auto_generated|divider|divider|op_5~3 ;
wire \Mod0|auto_generated|divider|divider|op_5~2_combout ;
wire \Mod0|auto_generated|divider|divider|op_5~5 ;
wire \Mod0|auto_generated|divider|divider|op_5~4_combout ;
wire \Mod0|auto_generated|divider|divider|op_5~7_cout ;
wire \Mod0|auto_generated|divider|divider|op_5~8_combout ;
wire \Mod1|auto_generated|divider|divider|op_2~1 ;
wire \Mod1|auto_generated|divider|divider|op_2~0_combout ;
wire \Mod1|auto_generated|divider|divider|op_2~3 ;
wire \Mod1|auto_generated|divider|divider|op_2~2_combout ;
wire \Mod1|auto_generated|divider|divider|op_2~5 ;
wire \Mod1|auto_generated|divider|divider|op_2~4_combout ;
wire \Mod1|auto_generated|divider|divider|op_2~7 ;
wire \Mod1|auto_generated|divider|divider|op_2~6_combout ;
wire \Mod1|auto_generated|divider|divider|op_2~8_combout ;
wire \integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ;
wire \integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ;
wire \stage_diff[1].auk_dsp_diff|dout_valid~q ;
wire \ena_diff_s[1]~0_combout ;
wire \stage_diff[0].auk_dsp_diff|dout_valid~q ;
wire \ena_diff_s[1]~q ;
wire \int_channel_cnt_inst|count[0]~q ;
wire \int_channel_cnt_inst|count[3]~q ;
wire \int_channel_cnt_inst|count[2]~q ;
wire \int_channel_cnt_inst|count[1]~q ;
wire \Mod2|auto_generated|divider|divider|StageOut[153]~0_combout ;
wire \Mod2|auto_generated|divider|divider|StageOut[153]~1_combout ;
wire \Mod2|auto_generated|divider|divider|StageOut[152]~2_combout ;
wire \Mod2|auto_generated|divider|divider|StageOut[152]~3_combout ;
wire \Mod2|auto_generated|divider|divider|StageOut[151]~4_combout ;
wire \Mod2|auto_generated|divider|divider|StageOut[151]~5_combout ;
wire \Mod2|auto_generated|divider|divider|StageOut[150]~6_combout ;
wire \Mod2|auto_generated|divider|divider|StageOut[150]~7_combout ;
wire \Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ;
wire \Mux18~0_combout ;
wire \Mux18~1_combout ;
wire \Mux18~2_combout ;
wire \Mux18~3_combout ;
wire \Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ;
wire \Mux18~4_combout ;
wire \Mux18~5_combout ;
wire \Mux18~6_combout ;
wire \Mux18~7_combout ;
wire \Mux18~8_combout ;
wire \Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ;
wire \Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ;
wire \Mux18~9_combout ;
wire \Mux0~0_combout ;
wire \Mux18~10_combout ;
wire \Mux17~2_combout ;
wire \Mux17~3_combout ;
wire \Mux17~4_combout ;
wire \Mux17~5_combout ;
wire \Mux17~6_combout ;
wire \Mux16~2_combout ;
wire \Mux16~3_combout ;
wire \Mux16~4_combout ;
wire \Mux16~5_combout ;
wire \Mux16~6_combout ;
wire \Mux15~2_combout ;
wire \Mux15~3_combout ;
wire \Mux15~4_combout ;
wire \Mux15~5_combout ;
wire \Mux15~6_combout ;
wire \Mux14~0_combout ;
wire \Mux14~1_combout ;
wire \Mux14~2_combout ;
wire \Mux14~3_combout ;
wire \Mux14~4_combout ;
wire \Mux14~5_combout ;
wire \Mux13~0_combout ;
wire \Mux13~1_combout ;
wire \Mux13~2_combout ;
wire \Mux13~3_combout ;
wire \Mux13~4_combout ;
wire \Mux13~5_combout ;
wire \Mux12~0_combout ;
wire \Mux12~1_combout ;
wire \Mux12~2_combout ;
wire \Mux12~3_combout ;
wire \Mux12~4_combout ;
wire \Mux12~5_combout ;
wire \Mux11~0_combout ;
wire \Mux11~1_combout ;
wire \Mux11~2_combout ;
wire \Mux11~3_combout ;
wire \Mux11~4_combout ;
wire \Mux11~5_combout ;
wire \Mux10~0_combout ;
wire \Mux10~1_combout ;
wire \Mux10~2_combout ;
wire \Mux10~3_combout ;
wire \Mux10~4_combout ;
wire \Mux10~5_combout ;
wire \Mux9~0_combout ;
wire \Mux9~1_combout ;
wire \Mux9~2_combout ;
wire \Mux9~3_combout ;
wire \Mux9~4_combout ;
wire \Mux9~5_combout ;
wire \Mux8~0_combout ;
wire \Mux8~1_combout ;
wire \Mux8~2_combout ;
wire \Mux8~3_combout ;
wire \Mux8~4_combout ;
wire \Mux8~5_combout ;
wire \Mux7~0_combout ;
wire \Mux7~1_combout ;
wire \Mux7~2_combout ;
wire \Mux7~3_combout ;
wire \Mux7~4_combout ;
wire \Mux7~5_combout ;
wire \Mux6~0_combout ;
wire \Mux6~1_combout ;
wire \Mux6~2_combout ;
wire \Mux6~3_combout ;
wire \Mux6~4_combout ;
wire \Mux6~5_combout ;
wire \Mux5~0_combout ;
wire \Mux5~1_combout ;
wire \Mux5~2_combout ;
wire \Mux5~3_combout ;
wire \Mux5~4_combout ;
wire \Mux5~5_combout ;
wire \Mux4~0_combout ;
wire \Mux4~1_combout ;
wire \Mux4~2_combout ;
wire \Mux4~3_combout ;
wire \Mux4~4_combout ;
wire \Mux4~5_combout ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \Mux3~2_combout ;
wire \Mux3~3_combout ;
wire \Mux3~4_combout ;
wire \Mux3~5_combout ;
wire \Mux2~0_combout ;
wire \Mux2~1_combout ;
wire \Mux2~2_combout ;
wire \Mux2~3_combout ;
wire \Mux2~4_combout ;
wire \Mux2~5_combout ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;
wire \Mux1~2_combout ;
wire \Mux1~3_combout ;
wire \Mux1~4_combout ;
wire \Mux1~5_combout ;
wire \Mux0~1_combout ;
wire \Mux0~2_combout ;
wire \Mux0~3_combout ;
wire \Mux0~4_combout ;
wire \Mux0~5_combout ;
wire \Mux0~6_combout ;
wire \ena_diff_s~1_combout ;
wire \ena_sample~0_combout ;
wire \integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~1_combout ;
wire \fifo_rdreq[5]~q ;
wire \fifo_rdreq[6]~q ;
wire \fifo_rdreq[4]~q ;
wire \fifo_rdreq[7]~q ;
wire \fifo_rdreq[2]~q ;
wire \fifo_rdreq[1]~q ;
wire \fifo_rdreq[0]~q ;
wire \fifo_rdreq[3]~q ;
wire \fifo_rdreq[8]~q ;
wire \ena_sample~1_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[10]~36_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[10]~37_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[9]~38_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[9]~39_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[8]~40_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[8]~41_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[14]~42_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[13]~43_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[12]~44_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[12]~45_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[18]~46_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[17]~47_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[16]~48_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[16]~49_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[20]~50_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[20]~51_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[21]~52_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[22]~53_combout ;
wire \ena_sample~2_combout ;
wire \ena_sample~3_combout ;
wire \ena_sample~4_combout ;
wire \ena_sample~5_combout ;
wire \sample_state~0_combout ;
wire \sample_state~1_combout ;
wire \Mod1|auto_generated|divider|divider|StageOut[12]~0_combout ;
wire \Mod1|auto_generated|divider|divider|StageOut[14]~1_combout ;
wire \always5~0_combout ;
wire \Mod1|auto_generated|divider|divider|StageOut[13]~2_combout ;
wire \always5~1_combout ;
wire \always5~2_combout ;
wire \always5~3_combout ;
wire \always5~4_combout ;
wire \always5~5_combout ;
wire \always5~6_combout ;
wire \always5~7_combout ;
wire \always5~8_combout ;
wire \always5~9_combout ;
wire \always5~10_combout ;
wire \Mux17~7_combout ;
wire \Mux16~7_combout ;
wire \Mux15~7_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[18]~54_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[22]~55_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[14]~56_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[13]~57_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[17]~58_combout ;
wire \Mod0|auto_generated|divider|divider|StageOut[21]~59_combout ;
wire \latency_cnt[3]~0_combout ;
wire \latency_cnt[0]~4_combout ;
wire \latency_cnt[0]~q ;
wire \latency_cnt[1]~3_combout ;
wire \latency_cnt[1]~q ;
wire \Add3~1_combout ;
wire \latency_cnt[2]~2_combout ;
wire \latency_cnt[2]~q ;
wire \Add3~0_combout ;
wire \latency_cnt[3]~1_combout ;
wire \latency_cnt[3]~q ;
wire \state~0_combout ;
wire \state~1_combout ;
wire \Add0~0_combout ;
wire \channel_out_int[1]~0_combout ;
wire \channel_out_int~1_combout ;
wire \channel_out_int[1]~2_combout ;
wire \channel_out_int~3_combout ;
wire \channel_out_int~4_combout ;
wire \Add0~1_combout ;
wire \channel_out_int~5_combout ;


cic_auk_dspip_integrator_14 \integrator[4].integrator_inner[2].integration (
	.register_fifofifo_data00(\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data001(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data019(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data021(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data031(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data041(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data051(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data061(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data071(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data081(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data091(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0101(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0111(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0121(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0131(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0141(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0151(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0181(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_13 \integrator[4].integrator_inner[1].integration (
	.register_fifofifo_data00(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[4].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data001(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data019(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data021(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data031(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data041(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data051(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data061(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data071(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data081(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data091(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0101(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0111(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0121(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0131(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0141(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0151(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0181(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_12 \integrator[4].integrator_inner[0].integration (
	.register_fifofifo_data00(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[4].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.q_b_4(q_b_4),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_channel_buffer_3 \integrator[3].fifo_regulator (
	.q({\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ,
\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ,\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ,
\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] }),
	.data({\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,
\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,
\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,
\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,
\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,
\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,
\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,
\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ,\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ,
\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ,\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ,
\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q }),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~1_combout ),
	.fifo_rdreq_3(\fifo_rdreq[3]~q ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_11 \integrator[3].integrator_inner[2].integration (
	.register_fifofifo_data00(\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[3].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data001(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data019(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data021(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data031(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data041(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data051(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data061(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data071(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data081(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data091(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0101(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0111(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0121(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0131(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0141(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0151(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0181(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_10 \integrator[3].integrator_inner[1].integration (
	.register_fifofifo_data00(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[3].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data001(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data019(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data021(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data031(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data041(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data051(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data061(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data071(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data081(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data091(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0101(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0111(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0121(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0131(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0141(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0151(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0181(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_9 \integrator[3].integrator_inner[0].integration (
	.register_fifofifo_data00(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[3].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.q_b_3(q_b_3),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_channel_buffer_2 \integrator[2].fifo_regulator (
	.q({\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ,
\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ,\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ,
\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] }),
	.data({\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,
\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,
\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,
\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,
\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,
\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,
\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,
\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ,\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ,
\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ,\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ,
\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q }),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~1_combout ),
	.fifo_rdreq_2(\fifo_rdreq[2]~q ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_8 \integrator[2].integrator_inner[2].integration (
	.register_fifofifo_data00(\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[2].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data001(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data019(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data021(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data031(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data041(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data051(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data061(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data071(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data081(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data091(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0101(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0111(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0121(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0131(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0141(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0151(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0181(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_7 \integrator[2].integrator_inner[1].integration (
	.register_fifofifo_data00(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[2].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data001(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data019(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data021(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data031(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data041(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data051(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data061(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data071(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data081(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data091(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0101(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0111(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0121(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0131(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0141(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0151(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0181(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_6 \integrator[2].integrator_inner[0].integration (
	.register_fifofifo_data00(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[2].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.q_b_2(q_b_2),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_channel_buffer_1 \integrator[1].fifo_regulator (
	.q({\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ,
\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ,\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ,
\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] }),
	.data({\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,
\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,
\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,
\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,
\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,
\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,
\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,
\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ,\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ,
\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ,\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ,
\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q }),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~1_combout ),
	.fifo_rdreq_1(\fifo_rdreq[1]~q ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_5 \integrator[1].integrator_inner[2].integration (
	.register_fifofifo_data00(\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[1].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data001(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data019(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data021(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data031(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data041(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data051(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data061(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data071(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data081(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data091(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0101(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0111(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0121(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0131(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0141(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0151(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0181(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_4 \integrator[1].integrator_inner[1].integration (
	.register_fifofifo_data00(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[1].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data001(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data019(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data021(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data031(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data041(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data051(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data061(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data071(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data081(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data091(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0101(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0111(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0121(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0131(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0141(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0151(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0181(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_3 \integrator[1].integrator_inner[0].integration (
	.register_fifofifo_data00(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[1].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.q_b_1(q_b_1),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_channel_buffer \integrator[0].fifo_regulator (
	.q({\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ,
\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ,\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ,
\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] }),
	.count_1(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[1]~q ),
	.count_2(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[2]~q ),
	.count_3(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[3]~q ),
	.count_4(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[4]~q ),
	.count_0(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[0]~q ),
	.count_5(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[5]~q ),
	.data({\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,
\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,
\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,
\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,
\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,
\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,
\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,
\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ,\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ,
\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ,\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ,
\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q }),
	.stall_reg(stall_reg),
	.ena_sample(\ena_sample~0_combout ),
	.valid_wreq(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~1_combout ),
	.fifo_rdreq_0(\fifo_rdreq[0]~q ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_downsample \integrator[0].j0.vrc_en_0.first_dsample (
	.sample_state_0(\sample_state[0]~q ),
	.count_6(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[6]~q ),
	.count_1(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[1]~q ),
	.count_2(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[2]~q ),
	.count_3(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[3]~q ),
	.count_4(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[4]~q ),
	.count_0(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[0]~q ),
	.count_5(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[5]~q ),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_2 \integrator[0].integrator_inner[2].integration (
	.register_fifofifo_data00(\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[0].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data001(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data019(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data021(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data031(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data041(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data051(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data061(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data071(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data081(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data091(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0101(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0111(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0121(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0131(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0141(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0151(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0181(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_1 \integrator[0].integrator_inner[1].integration (
	.register_fifofifo_data00(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[0].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data001(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data019(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data021(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data031(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data041(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data051(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data061(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data071(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data081(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data091(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0101(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0111(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0121(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0131(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0141(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0151(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0181(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator \integrator[0].integrator_inner[0].integration (
	.register_fifofifo_data00(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[0].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.q_b_0(q_b_0),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_differentiator_2 \stage_diff[2].auk_dsp_diff (
	.dout_0(dout_0),
	.dout_1(dout_1),
	.dout_2(dout_2),
	.dout_3(dout_3),
	.dout_4(dout_4),
	.dout_5(dout_5),
	.dout_6(dout_6),
	.dout_7(dout_7),
	.dout_8(dout_8),
	.dout_9(dout_9),
	.dout_10(dout_10),
	.dout_11(dout_11),
	.dout_12(dout_12),
	.dout_13(dout_13),
	.dout_14(dout_14),
	.dout_15(dout_15),
	.dout_16(dout_16),
	.dout_17(dout_17),
	.dout_18(dout_18),
	.dout_01(\stage_diff[1].auk_dsp_diff|dout[0]~q ),
	.dout_19(\stage_diff[1].auk_dsp_diff|dout[1]~q ),
	.dout_21(\stage_diff[1].auk_dsp_diff|dout[2]~q ),
	.dout_31(\stage_diff[1].auk_dsp_diff|dout[3]~q ),
	.dout_41(\stage_diff[1].auk_dsp_diff|dout[4]~q ),
	.dout_51(\stage_diff[1].auk_dsp_diff|dout[5]~q ),
	.dout_61(\stage_diff[1].auk_dsp_diff|dout[6]~q ),
	.dout_71(\stage_diff[1].auk_dsp_diff|dout[7]~q ),
	.dout_81(\stage_diff[1].auk_dsp_diff|dout[8]~q ),
	.dout_91(\stage_diff[1].auk_dsp_diff|dout[9]~q ),
	.dout_101(\stage_diff[1].auk_dsp_diff|dout[10]~q ),
	.dout_111(\stage_diff[1].auk_dsp_diff|dout[11]~q ),
	.dout_121(\stage_diff[1].auk_dsp_diff|dout[12]~q ),
	.dout_131(\stage_diff[1].auk_dsp_diff|dout[13]~q ),
	.dout_141(\stage_diff[1].auk_dsp_diff|dout[14]~q ),
	.dout_151(\stage_diff[1].auk_dsp_diff|dout[15]~q ),
	.dout_161(\stage_diff[1].auk_dsp_diff|dout[16]~q ),
	.dout_171(\stage_diff[1].auk_dsp_diff|dout[17]~q ),
	.dout_181(\stage_diff[1].auk_dsp_diff|dout[18]~q ),
	.stall_reg(stall_reg),
	.dout_valid1(dout_valid),
	.dout_valid2(\stage_diff[1].auk_dsp_diff|dout_valid~q ),
	.ena_diff_s_1(\ena_diff_s[1]~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_differentiator_1 \stage_diff[1].auk_dsp_diff (
	.dout_0(\stage_diff[1].auk_dsp_diff|dout[0]~q ),
	.dout_1(\stage_diff[1].auk_dsp_diff|dout[1]~q ),
	.dout_2(\stage_diff[1].auk_dsp_diff|dout[2]~q ),
	.dout_3(\stage_diff[1].auk_dsp_diff|dout[3]~q ),
	.dout_4(\stage_diff[1].auk_dsp_diff|dout[4]~q ),
	.dout_5(\stage_diff[1].auk_dsp_diff|dout[5]~q ),
	.dout_6(\stage_diff[1].auk_dsp_diff|dout[6]~q ),
	.dout_7(\stage_diff[1].auk_dsp_diff|dout[7]~q ),
	.dout_8(\stage_diff[1].auk_dsp_diff|dout[8]~q ),
	.dout_9(\stage_diff[1].auk_dsp_diff|dout[9]~q ),
	.dout_10(\stage_diff[1].auk_dsp_diff|dout[10]~q ),
	.dout_11(\stage_diff[1].auk_dsp_diff|dout[11]~q ),
	.dout_12(\stage_diff[1].auk_dsp_diff|dout[12]~q ),
	.dout_13(\stage_diff[1].auk_dsp_diff|dout[13]~q ),
	.dout_14(\stage_diff[1].auk_dsp_diff|dout[14]~q ),
	.dout_15(\stage_diff[1].auk_dsp_diff|dout[15]~q ),
	.dout_16(\stage_diff[1].auk_dsp_diff|dout[16]~q ),
	.dout_17(\stage_diff[1].auk_dsp_diff|dout[17]~q ),
	.dout_18(\stage_diff[1].auk_dsp_diff|dout[18]~q ),
	.dout_01(\stage_diff[0].auk_dsp_diff|dout[0]~q ),
	.dout_19(\stage_diff[0].auk_dsp_diff|dout[1]~q ),
	.dout_21(\stage_diff[0].auk_dsp_diff|dout[2]~q ),
	.dout_31(\stage_diff[0].auk_dsp_diff|dout[3]~q ),
	.dout_41(\stage_diff[0].auk_dsp_diff|dout[4]~q ),
	.dout_51(\stage_diff[0].auk_dsp_diff|dout[5]~q ),
	.dout_61(\stage_diff[0].auk_dsp_diff|dout[6]~q ),
	.dout_71(\stage_diff[0].auk_dsp_diff|dout[7]~q ),
	.dout_81(\stage_diff[0].auk_dsp_diff|dout[8]~q ),
	.dout_91(\stage_diff[0].auk_dsp_diff|dout[9]~q ),
	.dout_101(\stage_diff[0].auk_dsp_diff|dout[10]~q ),
	.dout_111(\stage_diff[0].auk_dsp_diff|dout[11]~q ),
	.dout_121(\stage_diff[0].auk_dsp_diff|dout[12]~q ),
	.dout_131(\stage_diff[0].auk_dsp_diff|dout[13]~q ),
	.dout_141(\stage_diff[0].auk_dsp_diff|dout[14]~q ),
	.dout_151(\stage_diff[0].auk_dsp_diff|dout[15]~q ),
	.dout_161(\stage_diff[0].auk_dsp_diff|dout[16]~q ),
	.dout_171(\stage_diff[0].auk_dsp_diff|dout[17]~q ),
	.dout_181(\stage_diff[0].auk_dsp_diff|dout[18]~q ),
	.stall_reg(stall_reg),
	.dout_valid1(\stage_diff[1].auk_dsp_diff|dout_valid~q ),
	.ena_diff_s_1(\ena_diff_s[1]~0_combout ),
	.dout_valid2(\stage_diff[0].auk_dsp_diff|dout_valid~q ),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_differentiator \stage_diff[0].auk_dsp_diff (
	.dout_0(\stage_diff[0].auk_dsp_diff|dout[0]~q ),
	.dout_1(\stage_diff[0].auk_dsp_diff|dout[1]~q ),
	.dout_2(\stage_diff[0].auk_dsp_diff|dout[2]~q ),
	.dout_3(\stage_diff[0].auk_dsp_diff|dout[3]~q ),
	.dout_4(\stage_diff[0].auk_dsp_diff|dout[4]~q ),
	.dout_5(\stage_diff[0].auk_dsp_diff|dout[5]~q ),
	.dout_6(\stage_diff[0].auk_dsp_diff|dout[6]~q ),
	.dout_7(\stage_diff[0].auk_dsp_diff|dout[7]~q ),
	.dout_8(\stage_diff[0].auk_dsp_diff|dout[8]~q ),
	.dout_9(\stage_diff[0].auk_dsp_diff|dout[9]~q ),
	.dout_10(\stage_diff[0].auk_dsp_diff|dout[10]~q ),
	.dout_11(\stage_diff[0].auk_dsp_diff|dout[11]~q ),
	.dout_12(\stage_diff[0].auk_dsp_diff|dout[12]~q ),
	.dout_13(\stage_diff[0].auk_dsp_diff|dout[13]~q ),
	.dout_14(\stage_diff[0].auk_dsp_diff|dout[14]~q ),
	.dout_15(\stage_diff[0].auk_dsp_diff|dout[15]~q ),
	.dout_16(\stage_diff[0].auk_dsp_diff|dout[16]~q ),
	.dout_17(\stage_diff[0].auk_dsp_diff|dout[17]~q ),
	.dout_18(\stage_diff[0].auk_dsp_diff|dout[18]~q ),
	.stall_reg(stall_reg),
	.ena_diff_s_1(\ena_diff_s[1]~0_combout ),
	.dout_valid1(\stage_diff[0].auk_dsp_diff|dout_valid~q ),
	.ena_diff_s_11(\ena_diff_s[1]~q ),
	.Mux18(\Mux18~10_combout ),
	.Mux14(\Mux14~5_combout ),
	.Mux13(\Mux13~5_combout ),
	.Mux12(\Mux12~5_combout ),
	.Mux11(\Mux11~5_combout ),
	.Mux10(\Mux10~5_combout ),
	.Mux9(\Mux9~5_combout ),
	.Mux8(\Mux8~5_combout ),
	.Mux7(\Mux7~5_combout ),
	.Mux6(\Mux6~5_combout ),
	.Mux5(\Mux5~5_combout ),
	.Mux4(\Mux4~5_combout ),
	.Mux3(\Mux3~5_combout ),
	.Mux2(\Mux2~5_combout ),
	.Mux1(\Mux1~5_combout ),
	.Mux0(\Mux0~6_combout ),
	.Mux17(\Mux17~7_combout ),
	.Mux16(\Mux16~7_combout ),
	.Mux15(\Mux15~7_combout ),
	.clk(clk),
	.reset_n(reset_n));

cic_counter_module_19 int_channel_cnt_inst(
	.ena_sample(\ena_sample~q ),
	.stall_reg(stall_reg),
	.count_0(\int_channel_cnt_inst|count[0]~q ),
	.count_3(\int_channel_cnt_inst|count[3]~q ),
	.count_2(\int_channel_cnt_inst|count[2]~q ),
	.count_1(\int_channel_cnt_inst|count[1]~q ),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_channel_buffer_8 \integrator[8].fifo_regulator (
	.q({\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ,
\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ,\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ,
\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] }),
	.data({\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,
\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,
\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,
\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,
\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,
\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,
\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,
\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ,\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ,
\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ,\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ,
\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q }),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~1_combout ),
	.fifo_rdreq_8(\fifo_rdreq[8]~q ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_26 \integrator[8].integrator_inner[2].integration (
	.register_fifofifo_data00(\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[8].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data001(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data019(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data021(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data031(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data041(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data051(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data061(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data071(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data081(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data091(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0101(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0111(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0121(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0131(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0141(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0151(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0181(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_25 \integrator[8].integrator_inner[1].integration (
	.register_fifofifo_data00(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[8].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data001(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data019(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data021(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data031(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data041(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data051(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data061(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data071(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data081(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data091(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0101(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0111(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0121(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0131(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0141(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0151(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0181(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_24 \integrator[8].integrator_inner[0].integration (
	.register_fifofifo_data00(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[8].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.q_b_8(q_b_8),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_channel_buffer_7 \integrator[7].fifo_regulator (
	.q({\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ,
\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ,\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ,
\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] }),
	.data({\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,
\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,
\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,
\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,
\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,
\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,
\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,
\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ,\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ,
\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ,\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ,
\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q }),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~1_combout ),
	.fifo_rdreq_7(\fifo_rdreq[7]~q ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_23 \integrator[7].integrator_inner[2].integration (
	.register_fifofifo_data00(\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[7].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data001(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data019(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data021(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data031(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data041(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data051(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data061(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data071(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data081(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data091(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0101(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0111(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0121(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0131(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0141(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0151(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0181(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_22 \integrator[7].integrator_inner[1].integration (
	.register_fifofifo_data00(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[7].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data001(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data019(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data021(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data031(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data041(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data051(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data061(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data071(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data081(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data091(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0101(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0111(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0121(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0131(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0141(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0151(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0181(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_21 \integrator[7].integrator_inner[0].integration (
	.register_fifofifo_data00(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[7].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.q_b_7(q_b_7),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_channel_buffer_6 \integrator[6].fifo_regulator (
	.q({\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ,
\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ,\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ,
\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] }),
	.data({\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,
\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,
\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,
\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,
\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,
\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,
\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,
\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ,\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ,
\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ,\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ,
\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q }),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~1_combout ),
	.fifo_rdreq_6(\fifo_rdreq[6]~q ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_20 \integrator[6].integrator_inner[2].integration (
	.register_fifofifo_data00(\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[6].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data001(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data019(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data021(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data031(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data041(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data051(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data061(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data071(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data081(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data091(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0101(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0111(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0121(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0131(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0141(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0151(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0181(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_19 \integrator[6].integrator_inner[1].integration (
	.register_fifofifo_data00(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[6].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data001(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data019(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data021(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data031(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data041(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data051(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data061(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data071(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data081(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data091(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0101(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0111(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0121(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0131(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0141(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0151(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0181(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_18 \integrator[6].integrator_inner[0].integration (
	.register_fifofifo_data00(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[6].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.q_b_6(q_b_6),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_channel_buffer_5 \integrator[5].fifo_regulator (
	.q({\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ,
\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ,\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ,
\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] }),
	.data({\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,
\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,
\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,
\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,
\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,
\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,
\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,
\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ,\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ,
\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ,\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ,
\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q }),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~1_combout ),
	.fifo_rdreq_5(\fifo_rdreq[5]~q ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_17 \integrator[5].integrator_inner[2].integration (
	.register_fifofifo_data00(\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[5].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data001(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data019(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data021(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data031(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data041(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data051(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data061(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data071(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data081(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data091(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0101(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0111(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0121(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0131(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0141(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0151(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0181(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_16 \integrator[5].integrator_inner[1].integration (
	.register_fifofifo_data00(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[5].integrator_inner[1].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.register_fifofifo_data001(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data019(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data021(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data031(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data041(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data051(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data061(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data071(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data081(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data091(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data0101(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data0111(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data0121(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data0131(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data0141(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data0151(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data0161(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data0171(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data0181(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_integrator_15 \integrator[5].integrator_inner[0].integration (
	.register_fifofifo_data00(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q ),
	.register_fifofifo_data01(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ),
	.register_fifofifo_data02(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ),
	.register_fifofifo_data03(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ),
	.register_fifofifo_data04(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ),
	.register_fifofifo_data05(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ),
	.register_fifofifo_data06(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ),
	.register_fifofifo_data07(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ),
	.register_fifofifo_data08(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ),
	.register_fifofifo_data09(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ),
	.register_fifofifo_data010(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ),
	.register_fifofifo_data011(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ),
	.register_fifofifo_data012(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ),
	.register_fifofifo_data013(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ),
	.register_fifofifo_data014(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ),
	.register_fifofifo_data015(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ),
	.register_fifofifo_data016(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ),
	.register_fifofifo_data017(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ),
	.register_fifofifo_data018(\integrator[5].integrator_inner[0].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ),
	.q_b_5(q_b_5),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

cic_auk_dspip_channel_buffer_4 \integrator[4].fifo_regulator (
	.q({\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ,
\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ,
\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ,
\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ,
\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ,
\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ,\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ,
\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] }),
	.data({\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][18]~q ,\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][17]~q ,
\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][16]~q ,\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][15]~q ,
\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][14]~q ,\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][13]~q ,
\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][12]~q ,\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][11]~q ,
\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][10]~q ,\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][9]~q ,
\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][8]~q ,\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][7]~q ,
\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][6]~q ,\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][5]~q ,
\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][4]~q ,\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][3]~q ,
\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][2]~q ,\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][1]~q ,
\integrator[4].integrator_inner[2].integration|glogic:integrator_pipeline_0_generate:u1|register_fifo:fifo_data[0][0]~q }),
	.stall_reg(stall_reg),
	.valid_wreq(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|valid_wreq~1_combout ),
	.fifo_rdreq_4(\fifo_rdreq[4]~q ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|op_24~0 (
	.dataa(\int_channel_cnt_inst|count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Mod2|auto_generated|divider|divider|op_24~0_combout ),
	.cout(\Mod2|auto_generated|divider|divider|op_24~1 ));
defparam \Mod2|auto_generated|divider|divider|op_24~0 .lut_mask = 16'h55AA;
defparam \Mod2|auto_generated|divider|divider|op_24~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|op_23~0 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Mod2|auto_generated|divider|divider|op_23~0_combout ),
	.cout(\Mod2|auto_generated|divider|divider|op_23~1 ));
defparam \Mod2|auto_generated|divider|divider|op_23~0 .lut_mask = 16'h55AA;
defparam \Mod2|auto_generated|divider|divider|op_23~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|op_23~2 (
	.dataa(\int_channel_cnt_inst|count[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod2|auto_generated|divider|divider|op_23~1 ),
	.combout(\Mod2|auto_generated|divider|divider|op_23~2_combout ),
	.cout(\Mod2|auto_generated|divider|divider|op_23~3 ));
defparam \Mod2|auto_generated|divider|divider|op_23~2 .lut_mask = 16'h5A5F;
defparam \Mod2|auto_generated|divider|divider|op_23~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|op_23~4 (
	.dataa(\int_channel_cnt_inst|count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod2|auto_generated|divider|divider|op_23~3 ),
	.combout(\Mod2|auto_generated|divider|divider|op_23~4_combout ),
	.cout(\Mod2|auto_generated|divider|divider|op_23~5 ));
defparam \Mod2|auto_generated|divider|divider|op_23~4 .lut_mask = 16'h5A5F;
defparam \Mod2|auto_generated|divider|divider|op_23~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|op_23~6 (
	.dataa(\int_channel_cnt_inst|count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod2|auto_generated|divider|divider|op_23~5 ),
	.combout(\Mod2|auto_generated|divider|divider|op_23~6_combout ),
	.cout(\Mod2|auto_generated|divider|divider|op_23~7 ));
defparam \Mod2|auto_generated|divider|divider|op_23~6 .lut_mask = 16'h5A5F;
defparam \Mod2|auto_generated|divider|divider|op_23~6 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|op_23~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod2|auto_generated|divider|divider|op_23~7 ),
	.combout(),
	.cout(\Mod2|auto_generated|divider|divider|op_23~9_cout ));
defparam \Mod2|auto_generated|divider|divider|op_23~9 .lut_mask = 16'h000F;
defparam \Mod2|auto_generated|divider|divider|op_23~9 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|op_23~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Mod2|auto_generated|divider|divider|op_23~9_cout ),
	.combout(\Mod2|auto_generated|divider|divider|op_23~10_combout ),
	.cout());
defparam \Mod2|auto_generated|divider|divider|op_23~10 .lut_mask = 16'h0F0F;
defparam \Mod2|auto_generated|divider|divider|op_23~10 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|op_24~2 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[150]~6_combout ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[150]~7_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod2|auto_generated|divider|divider|op_24~1 ),
	.combout(\Mod2|auto_generated|divider|divider|op_24~2_combout ),
	.cout(\Mod2|auto_generated|divider|divider|op_24~3 ));
defparam \Mod2|auto_generated|divider|divider|op_24~2 .lut_mask = 16'h967F;
defparam \Mod2|auto_generated|divider|divider|op_24~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|op_24~4 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[151]~4_combout ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[151]~5_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod2|auto_generated|divider|divider|op_24~3 ),
	.combout(\Mod2|auto_generated|divider|divider|op_24~4_combout ),
	.cout(\Mod2|auto_generated|divider|divider|op_24~5 ));
defparam \Mod2|auto_generated|divider|divider|op_24~4 .lut_mask = 16'h96EF;
defparam \Mod2|auto_generated|divider|divider|op_24~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|op_24~6 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[152]~2_combout ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[152]~3_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod2|auto_generated|divider|divider|op_24~5 ),
	.combout(\Mod2|auto_generated|divider|divider|op_24~6_combout ),
	.cout(\Mod2|auto_generated|divider|divider|op_24~7 ));
defparam \Mod2|auto_generated|divider|divider|op_24~6 .lut_mask = 16'h967F;
defparam \Mod2|auto_generated|divider|divider|op_24~6 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|op_24~9 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[153]~0_combout ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[153]~1_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod2|auto_generated|divider|divider|op_24~7 ),
	.combout(),
	.cout(\Mod2|auto_generated|divider|divider|op_24~9_cout ));
defparam \Mod2|auto_generated|divider|divider|op_24~9 .lut_mask = 16'h00EF;
defparam \Mod2|auto_generated|divider|divider|op_24~9 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|op_24~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Mod2|auto_generated|divider|divider|op_24~9_cout ),
	.combout(\Mod2|auto_generated|divider|divider|op_24~10_combout ),
	.cout());
defparam \Mod2|auto_generated|divider|divider|op_24~10 .lut_mask = 16'h0F0F;
defparam \Mod2|auto_generated|divider|divider|op_24~10 .sum_lutc_input = "cin";

dffeas ena_sample(
	.clk(clk),
	.d(\ena_sample~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\ena_sample~q ),
	.prn(vcc));
defparam ena_sample.is_wysiwyg = "true";
defparam ena_sample.power_up = "low";

dffeas \sample_state[0] (
	.clk(clk),
	.d(\sample_state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\sample_state[0]~q ),
	.prn(vcc));
defparam \sample_state[0] .is_wysiwyg = "true";
defparam \sample_state[0] .power_up = "low";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_5~0 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|op_5~0_combout ),
	.cout(\Mod0|auto_generated|divider|divider|op_5~1 ));
defparam \Mod0|auto_generated|divider|divider|op_5~0 .lut_mask = 16'h55AA;
defparam \Mod0|auto_generated|divider|divider|op_5~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_1~0 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|op_1~0_combout ),
	.cout(\Mod0|auto_generated|divider|divider|op_1~1 ));
defparam \Mod0|auto_generated|divider|divider|op_1~0 .lut_mask = 16'h55AA;
defparam \Mod0|auto_generated|divider|divider|op_1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_1~2 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|op_1~1 ),
	.combout(\Mod0|auto_generated|divider|divider|op_1~2_combout ),
	.cout(\Mod0|auto_generated|divider|divider|op_1~3 ));
defparam \Mod0|auto_generated|divider|divider|op_1~2 .lut_mask = 16'h5A5F;
defparam \Mod0|auto_generated|divider|divider|op_1~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_1~4 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|op_1~3 ),
	.combout(\Mod0|auto_generated|divider|divider|op_1~4_combout ),
	.cout(\Mod0|auto_generated|divider|divider|op_1~5 ));
defparam \Mod0|auto_generated|divider|divider|op_1~4 .lut_mask = 16'h5AAF;
defparam \Mod0|auto_generated|divider|divider|op_1~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_1~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Mod0|auto_generated|divider|divider|op_1~5 ),
	.combout(\Mod0|auto_generated|divider|divider|op_1~6_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|op_1~6 .lut_mask = 16'h0F0F;
defparam \Mod0|auto_generated|divider|divider|op_1~6 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_2~0 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|op_2~0_combout ),
	.cout(\Mod0|auto_generated|divider|divider|op_2~1 ));
defparam \Mod0|auto_generated|divider|divider|op_2~0 .lut_mask = 16'h55AA;
defparam \Mod0|auto_generated|divider|divider|op_2~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_2~2 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[8]~40_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[8]~41_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|op_2~1 ),
	.combout(\Mod0|auto_generated|divider|divider|op_2~2_combout ),
	.cout(\Mod0|auto_generated|divider|divider|op_2~3 ));
defparam \Mod0|auto_generated|divider|divider|op_2~2 .lut_mask = 16'h967F;
defparam \Mod0|auto_generated|divider|divider|op_2~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_2~4 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[9]~38_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[9]~39_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|op_2~3 ),
	.combout(\Mod0|auto_generated|divider|divider|op_2~4_combout ),
	.cout(\Mod0|auto_generated|divider|divider|op_2~5 ));
defparam \Mod0|auto_generated|divider|divider|op_2~4 .lut_mask = 16'h96EF;
defparam \Mod0|auto_generated|divider|divider|op_2~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_2~7 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[10]~36_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[10]~37_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|op_2~5 ),
	.combout(),
	.cout(\Mod0|auto_generated|divider|divider|op_2~7_cout ));
defparam \Mod0|auto_generated|divider|divider|op_2~7 .lut_mask = 16'h007F;
defparam \Mod0|auto_generated|divider|divider|op_2~7 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_2~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Mod0|auto_generated|divider|divider|op_2~7_cout ),
	.combout(\Mod0|auto_generated|divider|divider|op_2~8_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|op_2~8 .lut_mask = 16'hF0F0;
defparam \Mod0|auto_generated|divider|divider|op_2~8 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_3~0 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|op_3~0_combout ),
	.cout(\Mod0|auto_generated|divider|divider|op_3~1 ));
defparam \Mod0|auto_generated|divider|divider|op_3~0 .lut_mask = 16'h55AA;
defparam \Mod0|auto_generated|divider|divider|op_3~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_3~2 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[12]~44_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[12]~45_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|op_3~1 ),
	.combout(\Mod0|auto_generated|divider|divider|op_3~2_combout ),
	.cout(\Mod0|auto_generated|divider|divider|op_3~3 ));
defparam \Mod0|auto_generated|divider|divider|op_3~2 .lut_mask = 16'h967F;
defparam \Mod0|auto_generated|divider|divider|op_3~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_3~4 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[13]~57_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[13]~43_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|op_3~3 ),
	.combout(\Mod0|auto_generated|divider|divider|op_3~4_combout ),
	.cout(\Mod0|auto_generated|divider|divider|op_3~5 ));
defparam \Mod0|auto_generated|divider|divider|op_3~4 .lut_mask = 16'h96EF;
defparam \Mod0|auto_generated|divider|divider|op_3~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_3~7 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[14]~56_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[14]~42_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|op_3~5 ),
	.combout(),
	.cout(\Mod0|auto_generated|divider|divider|op_3~7_cout ));
defparam \Mod0|auto_generated|divider|divider|op_3~7 .lut_mask = 16'h007F;
defparam \Mod0|auto_generated|divider|divider|op_3~7 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_3~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Mod0|auto_generated|divider|divider|op_3~7_cout ),
	.combout(\Mod0|auto_generated|divider|divider|op_3~8_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|op_3~8 .lut_mask = 16'hF0F0;
defparam \Mod0|auto_generated|divider|divider|op_3~8 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_4~0 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|op_4~0_combout ),
	.cout(\Mod0|auto_generated|divider|divider|op_4~1 ));
defparam \Mod0|auto_generated|divider|divider|op_4~0 .lut_mask = 16'h55AA;
defparam \Mod0|auto_generated|divider|divider|op_4~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_4~2 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[16]~48_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[16]~49_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|op_4~1 ),
	.combout(\Mod0|auto_generated|divider|divider|op_4~2_combout ),
	.cout(\Mod0|auto_generated|divider|divider|op_4~3 ));
defparam \Mod0|auto_generated|divider|divider|op_4~2 .lut_mask = 16'h967F;
defparam \Mod0|auto_generated|divider|divider|op_4~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_4~4 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[17]~58_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[17]~47_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|op_4~3 ),
	.combout(\Mod0|auto_generated|divider|divider|op_4~4_combout ),
	.cout(\Mod0|auto_generated|divider|divider|op_4~5 ));
defparam \Mod0|auto_generated|divider|divider|op_4~4 .lut_mask = 16'h96EF;
defparam \Mod0|auto_generated|divider|divider|op_4~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_4~7 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[18]~54_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[18]~46_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|op_4~5 ),
	.combout(),
	.cout(\Mod0|auto_generated|divider|divider|op_4~7_cout ));
defparam \Mod0|auto_generated|divider|divider|op_4~7 .lut_mask = 16'h007F;
defparam \Mod0|auto_generated|divider|divider|op_4~7 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_4~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Mod0|auto_generated|divider|divider|op_4~7_cout ),
	.combout(\Mod0|auto_generated|divider|divider|op_4~8_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|op_4~8 .lut_mask = 16'hF0F0;
defparam \Mod0|auto_generated|divider|divider|op_4~8 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_5~2 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[20]~50_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[20]~51_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|op_5~1 ),
	.combout(\Mod0|auto_generated|divider|divider|op_5~2_combout ),
	.cout(\Mod0|auto_generated|divider|divider|op_5~3 ));
defparam \Mod0|auto_generated|divider|divider|op_5~2 .lut_mask = 16'h967F;
defparam \Mod0|auto_generated|divider|divider|op_5~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_5~4 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[21]~59_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[21]~52_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|op_5~3 ),
	.combout(\Mod0|auto_generated|divider|divider|op_5~4_combout ),
	.cout(\Mod0|auto_generated|divider|divider|op_5~5 ));
defparam \Mod0|auto_generated|divider|divider|op_5~4 .lut_mask = 16'h96EF;
defparam \Mod0|auto_generated|divider|divider|op_5~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_5~7 (
	.dataa(\Mod0|auto_generated|divider|divider|StageOut[22]~55_combout ),
	.datab(\Mod0|auto_generated|divider|divider|StageOut[22]~53_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod0|auto_generated|divider|divider|op_5~5 ),
	.combout(),
	.cout(\Mod0|auto_generated|divider|divider|op_5~7_cout ));
defparam \Mod0|auto_generated|divider|divider|op_5~7 .lut_mask = 16'h007F;
defparam \Mod0|auto_generated|divider|divider|op_5~7 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|op_5~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Mod0|auto_generated|divider|divider|op_5~7_cout ),
	.combout(\Mod0|auto_generated|divider|divider|op_5~8_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|op_5~8 .lut_mask = 16'hF0F0;
defparam \Mod0|auto_generated|divider|divider|op_5~8 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod1|auto_generated|divider|divider|op_2~0 (
	.dataa(\int_channel_cnt_inst|count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Mod1|auto_generated|divider|divider|op_2~0_combout ),
	.cout(\Mod1|auto_generated|divider|divider|op_2~1 ));
defparam \Mod1|auto_generated|divider|divider|op_2~0 .lut_mask = 16'h55AA;
defparam \Mod1|auto_generated|divider|divider|op_2~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod1|auto_generated|divider|divider|op_2~2 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod1|auto_generated|divider|divider|op_2~1 ),
	.combout(\Mod1|auto_generated|divider|divider|op_2~2_combout ),
	.cout(\Mod1|auto_generated|divider|divider|op_2~3 ));
defparam \Mod1|auto_generated|divider|divider|op_2~2 .lut_mask = 16'h5A5F;
defparam \Mod1|auto_generated|divider|divider|op_2~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod1|auto_generated|divider|divider|op_2~4 (
	.dataa(\int_channel_cnt_inst|count[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod1|auto_generated|divider|divider|op_2~3 ),
	.combout(\Mod1|auto_generated|divider|divider|op_2~4_combout ),
	.cout(\Mod1|auto_generated|divider|divider|op_2~5 ));
defparam \Mod1|auto_generated|divider|divider|op_2~4 .lut_mask = 16'h5AAF;
defparam \Mod1|auto_generated|divider|divider|op_2~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod1|auto_generated|divider|divider|op_2~6 (
	.dataa(\int_channel_cnt_inst|count[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Mod1|auto_generated|divider|divider|op_2~5 ),
	.combout(\Mod1|auto_generated|divider|divider|op_2~6_combout ),
	.cout(\Mod1|auto_generated|divider|divider|op_2~7 ));
defparam \Mod1|auto_generated|divider|divider|op_2~6 .lut_mask = 16'h5A5F;
defparam \Mod1|auto_generated|divider|divider|op_2~6 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Mod1|auto_generated|divider|divider|op_2~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Mod1|auto_generated|divider|divider|op_2~7 ),
	.combout(\Mod1|auto_generated|divider|divider|op_2~8_combout ),
	.cout());
defparam \Mod1|auto_generated|divider|divider|op_2~8 .lut_mask = 16'hF0F0;
defparam \Mod1|auto_generated|divider|divider|op_2~8 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \ena_diff_s[1]~0 (
	.dataa(reset_n),
	.datab(stall_reg),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ena_diff_s[1]~0_combout ),
	.cout());
defparam \ena_diff_s[1]~0 .lut_mask = 16'h7777;
defparam \ena_diff_s[1]~0 .sum_lutc_input = "datac";

dffeas \ena_diff_s[1] (
	.clk(clk),
	.d(\ena_diff_s~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ena_diff_s[1]~0_combout ),
	.q(\ena_diff_s[1]~q ),
	.prn(vcc));
defparam \ena_diff_s[1] .is_wysiwyg = "true";
defparam \ena_diff_s[1] .power_up = "low";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|StageOut[153]~0 (
	.dataa(\int_channel_cnt_inst|count[3]~q ),
	.datab(\Mod2|auto_generated|divider|divider|op_23~10_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mod2|auto_generated|divider|divider|StageOut[153]~0_combout ),
	.cout());
defparam \Mod2|auto_generated|divider|divider|StageOut[153]~0 .lut_mask = 16'hEEEE;
defparam \Mod2|auto_generated|divider|divider|StageOut[153]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|StageOut[153]~1 (
	.dataa(\Mod2|auto_generated|divider|divider|op_23~6_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod2|auto_generated|divider|divider|op_23~10_combout ),
	.cin(gnd),
	.combout(\Mod2|auto_generated|divider|divider|StageOut[153]~1_combout ),
	.cout());
defparam \Mod2|auto_generated|divider|divider|StageOut[153]~1 .lut_mask = 16'hAAFF;
defparam \Mod2|auto_generated|divider|divider|StageOut[153]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|StageOut[152]~2 (
	.dataa(\Mod2|auto_generated|divider|divider|op_23~10_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\int_channel_cnt_inst|count[3]~q ),
	.cin(gnd),
	.combout(\Mod2|auto_generated|divider|divider|StageOut[152]~2_combout ),
	.cout());
defparam \Mod2|auto_generated|divider|divider|StageOut[152]~2 .lut_mask = 16'hAAFF;
defparam \Mod2|auto_generated|divider|divider|StageOut[152]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|StageOut[152]~3 (
	.dataa(\Mod2|auto_generated|divider|divider|op_23~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod2|auto_generated|divider|divider|op_23~10_combout ),
	.cin(gnd),
	.combout(\Mod2|auto_generated|divider|divider|StageOut[152]~3_combout ),
	.cout());
defparam \Mod2|auto_generated|divider|divider|StageOut[152]~3 .lut_mask = 16'hAAFF;
defparam \Mod2|auto_generated|divider|divider|StageOut[152]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|StageOut[151]~4 (
	.dataa(\int_channel_cnt_inst|count[2]~q ),
	.datab(\Mod2|auto_generated|divider|divider|op_23~10_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mod2|auto_generated|divider|divider|StageOut[151]~4_combout ),
	.cout());
defparam \Mod2|auto_generated|divider|divider|StageOut[151]~4 .lut_mask = 16'hEEEE;
defparam \Mod2|auto_generated|divider|divider|StageOut[151]~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|StageOut[151]~5 (
	.dataa(\Mod2|auto_generated|divider|divider|op_23~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod2|auto_generated|divider|divider|op_23~10_combout ),
	.cin(gnd),
	.combout(\Mod2|auto_generated|divider|divider|StageOut[151]~5_combout ),
	.cout());
defparam \Mod2|auto_generated|divider|divider|StageOut[151]~5 .lut_mask = 16'hAAFF;
defparam \Mod2|auto_generated|divider|divider|StageOut[151]~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|StageOut[150]~6 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\Mod2|auto_generated|divider|divider|op_23~10_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mod2|auto_generated|divider|divider|StageOut[150]~6_combout ),
	.cout());
defparam \Mod2|auto_generated|divider|divider|StageOut[150]~6 .lut_mask = 16'hEEEE;
defparam \Mod2|auto_generated|divider|divider|StageOut[150]~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|StageOut[150]~7 (
	.dataa(\Mod2|auto_generated|divider|divider|op_23~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod2|auto_generated|divider|divider|op_23~10_combout ),
	.cin(gnd),
	.combout(\Mod2|auto_generated|divider|divider|StageOut[150]~7_combout ),
	.cout());
defparam \Mod2|auto_generated|divider|divider|StageOut[150]~7 .lut_mask = 16'hAAFF;
defparam \Mod2|auto_generated|divider|divider|StageOut[150]~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|StageOut[155]~8 (
	.dataa(\int_channel_cnt_inst|count[0]~q ),
	.datab(\Mod2|auto_generated|divider|divider|op_24~0_combout ),
	.datac(gnd),
	.datad(\Mod2|auto_generated|divider|divider|op_24~10_combout ),
	.cin(gnd),
	.combout(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.cout());
defparam \Mod2|auto_generated|divider|divider|StageOut[155]~8 .lut_mask = 16'hAACC;
defparam \Mod2|auto_generated|divider|divider|StageOut[155]~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux18~0 (
	.dataa(\int_channel_cnt_inst|count[0]~q ),
	.datab(\Mod2|auto_generated|divider|divider|op_24~0_combout ),
	.datac(\Mod2|auto_generated|divider|divider|op_24~10_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux18~0_combout ),
	.cout());
defparam \Mux18~0 .lut_mask = 16'hACAC;
defparam \Mux18~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux18~1 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[150]~6_combout ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[150]~7_combout ),
	.datac(\Mod2|auto_generated|divider|divider|op_24~2_combout ),
	.datad(\Mod2|auto_generated|divider|divider|op_24~10_combout ),
	.cin(gnd),
	.combout(\Mux18~1_combout ),
	.cout());
defparam \Mux18~1 .lut_mask = 16'hFAFC;
defparam \Mux18~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux18~2 (
	.dataa(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datab(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datac(\Mux18~0_combout ),
	.datad(\Mux18~1_combout ),
	.cin(gnd),
	.combout(\Mux18~2_combout ),
	.cout());
defparam \Mux18~2 .lut_mask = 16'hEFFE;
defparam \Mux18~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux18~3 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datac(\Mux18~2_combout ),
	.datad(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.cin(gnd),
	.combout(\Mux18~3_combout ),
	.cout());
defparam \Mux18~3 .lut_mask = 16'hFFBE;
defparam \Mux18~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|StageOut[156]~9 (
	.dataa(\Mod2|auto_generated|divider|divider|op_24~2_combout ),
	.datab(\Mod2|auto_generated|divider|divider|op_24~10_combout ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[150]~6_combout ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[150]~7_combout ),
	.cin(gnd),
	.combout(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.cout());
defparam \Mod2|auto_generated|divider|divider|StageOut[156]~9 .lut_mask = 16'hFFB8;
defparam \Mod2|auto_generated|divider|divider|StageOut[156]~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux18~4 (
	.dataa(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[150]~6_combout ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[150]~7_combout ),
	.datad(\int_channel_cnt_inst|count[0]~q ),
	.cin(gnd),
	.combout(\Mux18~4_combout ),
	.cout());
defparam \Mux18~4 .lut_mask = 16'hEBBE;
defparam \Mux18~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux18~5 (
	.dataa(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datab(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datac(\Mod2|auto_generated|divider|divider|op_24~2_combout ),
	.datad(\Mod2|auto_generated|divider|divider|op_24~0_combout ),
	.cin(gnd),
	.combout(\Mux18~5_combout ),
	.cout());
defparam \Mux18~5 .lut_mask = 16'hEFFE;
defparam \Mux18~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux18~6 (
	.dataa(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datab(\int_channel_cnt_inst|count[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux18~6_combout ),
	.cout());
defparam \Mux18~6 .lut_mask = 16'hEEEE;
defparam \Mux18~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux18~7 (
	.dataa(\Mod2|auto_generated|divider|divider|op_24~10_combout ),
	.datab(\Mux18~4_combout ),
	.datac(\Mux18~5_combout ),
	.datad(\Mux18~6_combout ),
	.cin(gnd),
	.combout(\Mux18~7_combout ),
	.cout());
defparam \Mux18~7 .lut_mask = 16'hFFD8;
defparam \Mux18~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux18~8 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datac(\Mux18~7_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.cin(gnd),
	.combout(\Mux18~8_combout ),
	.cout());
defparam \Mux18~8 .lut_mask = 16'hFFBE;
defparam \Mux18~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|StageOut[157]~10 (
	.dataa(\Mod2|auto_generated|divider|divider|op_24~4_combout ),
	.datab(\Mod2|auto_generated|divider|divider|op_24~10_combout ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[151]~4_combout ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[151]~5_combout ),
	.cin(gnd),
	.combout(\Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ),
	.cout());
defparam \Mod2|auto_generated|divider|divider|StageOut[157]~10 .lut_mask = 16'hFFB8;
defparam \Mod2|auto_generated|divider|divider|StageOut[157]~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod2|auto_generated|divider|divider|StageOut[158]~11 (
	.dataa(\Mod2|auto_generated|divider|divider|op_24~6_combout ),
	.datab(\Mod2|auto_generated|divider|divider|op_24~10_combout ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[152]~2_combout ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[152]~3_combout ),
	.cin(gnd),
	.combout(\Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ),
	.cout());
defparam \Mod2|auto_generated|divider|divider|StageOut[158]~11 .lut_mask = 16'hFFB8;
defparam \Mod2|auto_generated|divider|divider|StageOut[158]~11 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux18~9 (
	.dataa(\Mux18~3_combout ),
	.datab(\Mux18~8_combout ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ),
	.cin(gnd),
	.combout(\Mux18~9_combout ),
	.cout());
defparam \Mux18~9 .lut_mask = 16'hACFF;
defparam \Mux18~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux0~0 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hBFFF;
defparam \Mux0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux18~10 (
	.dataa(\Mux18~9_combout ),
	.datab(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.datac(\Mux0~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux18~10_combout ),
	.cout());
defparam \Mux18~10 .lut_mask = 16'hFEFE;
defparam \Mux18~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux17~2 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datab(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datac(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.cin(gnd),
	.combout(\Mux17~2_combout ),
	.cout());
defparam \Mux17~2 .lut_mask = 16'hFDFE;
defparam \Mux17~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux17~3 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datab(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datad(\Mux17~2_combout ),
	.cin(gnd),
	.combout(\Mux17~3_combout ),
	.cout());
defparam \Mux17~3 .lut_mask = 16'hEFFE;
defparam \Mux17~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux17~4 (
	.dataa(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datac(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.cin(gnd),
	.combout(\Mux17~4_combout ),
	.cout());
defparam \Mux17~4 .lut_mask = 16'hFBFE;
defparam \Mux17~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux17~5 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datab(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datad(\Mux17~4_combout ),
	.cin(gnd),
	.combout(\Mux17~5_combout ),
	.cout());
defparam \Mux17~5 .lut_mask = 16'hEFFE;
defparam \Mux17~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux17~6 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ),
	.datab(\Mux17~3_combout ),
	.datac(\Mux17~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux17~6_combout ),
	.cout());
defparam \Mux17~6 .lut_mask = 16'hD8D8;
defparam \Mux17~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux16~2 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datab(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datac(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.cin(gnd),
	.combout(\Mux16~2_combout ),
	.cout());
defparam \Mux16~2 .lut_mask = 16'hFDFE;
defparam \Mux16~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux16~3 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datab(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datad(\Mux16~2_combout ),
	.cin(gnd),
	.combout(\Mux16~3_combout ),
	.cout());
defparam \Mux16~3 .lut_mask = 16'hEFFE;
defparam \Mux16~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux16~4 (
	.dataa(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datac(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.cin(gnd),
	.combout(\Mux16~4_combout ),
	.cout());
defparam \Mux16~4 .lut_mask = 16'hFBFE;
defparam \Mux16~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux16~5 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datab(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datad(\Mux16~4_combout ),
	.cin(gnd),
	.combout(\Mux16~5_combout ),
	.cout());
defparam \Mux16~5 .lut_mask = 16'hEFFE;
defparam \Mux16~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux16~6 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ),
	.datab(\Mux16~3_combout ),
	.datac(\Mux16~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux16~6_combout ),
	.cout());
defparam \Mux16~6 .lut_mask = 16'hD8D8;
defparam \Mux16~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux15~2 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datab(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datac(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.cin(gnd),
	.combout(\Mux15~2_combout ),
	.cout());
defparam \Mux15~2 .lut_mask = 16'hFDFE;
defparam \Mux15~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux15~3 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datab(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datad(\Mux15~2_combout ),
	.cin(gnd),
	.combout(\Mux15~3_combout ),
	.cout());
defparam \Mux15~3 .lut_mask = 16'hEFFE;
defparam \Mux15~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux15~4 (
	.dataa(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datac(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.cin(gnd),
	.combout(\Mux15~4_combout ),
	.cout());
defparam \Mux15~4 .lut_mask = 16'hFBFE;
defparam \Mux15~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux15~5 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datab(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datad(\Mux15~4_combout ),
	.cin(gnd),
	.combout(\Mux15~5_combout ),
	.cout());
defparam \Mux15~5 .lut_mask = 16'hEFFE;
defparam \Mux15~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux15~6 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ),
	.datab(\Mux15~3_combout ),
	.datac(\Mux15~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux15~6_combout ),
	.cout());
defparam \Mux15~6 .lut_mask = 16'hD8D8;
defparam \Mux15~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux14~0 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datab(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.cin(gnd),
	.combout(\Mux14~0_combout ),
	.cout());
defparam \Mux14~0 .lut_mask = 16'hFFDE;
defparam \Mux14~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux14~1 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datac(\Mux14~0_combout ),
	.datad(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.cin(gnd),
	.combout(\Mux14~1_combout ),
	.cout());
defparam \Mux14~1 .lut_mask = 16'hFFBE;
defparam \Mux14~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux14~2 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datab(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.cin(gnd),
	.combout(\Mux14~2_combout ),
	.cout());
defparam \Mux14~2 .lut_mask = 16'hFFDE;
defparam \Mux14~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux14~3 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datac(\Mux14~2_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.cin(gnd),
	.combout(\Mux14~3_combout ),
	.cout());
defparam \Mux14~3 .lut_mask = 16'hFFBE;
defparam \Mux14~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux14~4 (
	.dataa(\Mux14~1_combout ),
	.datab(\Mux14~3_combout ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ),
	.cin(gnd),
	.combout(\Mux14~4_combout ),
	.cout());
defparam \Mux14~4 .lut_mask = 16'hACFF;
defparam \Mux14~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux14~5 (
	.dataa(\Mux14~4_combout ),
	.datab(\Mux0~0_combout ),
	.datac(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux14~5_combout ),
	.cout());
defparam \Mux14~5 .lut_mask = 16'hFEFE;
defparam \Mux14~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux13~0 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datab(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
defparam \Mux13~0 .lut_mask = 16'hFFDE;
defparam \Mux13~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux13~1 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datac(\Mux13~0_combout ),
	.datad(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.cin(gnd),
	.combout(\Mux13~1_combout ),
	.cout());
defparam \Mux13~1 .lut_mask = 16'hFFBE;
defparam \Mux13~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux13~2 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datab(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.cin(gnd),
	.combout(\Mux13~2_combout ),
	.cout());
defparam \Mux13~2 .lut_mask = 16'hFFDE;
defparam \Mux13~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux13~3 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datac(\Mux13~2_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.cin(gnd),
	.combout(\Mux13~3_combout ),
	.cout());
defparam \Mux13~3 .lut_mask = 16'hFFBE;
defparam \Mux13~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux13~4 (
	.dataa(\Mux13~1_combout ),
	.datab(\Mux13~3_combout ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ),
	.cin(gnd),
	.combout(\Mux13~4_combout ),
	.cout());
defparam \Mux13~4 .lut_mask = 16'hACFF;
defparam \Mux13~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux13~5 (
	.dataa(\Mux13~4_combout ),
	.datab(\Mux0~0_combout ),
	.datac(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux13~5_combout ),
	.cout());
defparam \Mux13~5 .lut_mask = 16'hFEFE;
defparam \Mux13~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux12~0 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datab(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
defparam \Mux12~0 .lut_mask = 16'hFFDE;
defparam \Mux12~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux12~1 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datac(\Mux12~0_combout ),
	.datad(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.cin(gnd),
	.combout(\Mux12~1_combout ),
	.cout());
defparam \Mux12~1 .lut_mask = 16'hFFBE;
defparam \Mux12~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux12~2 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datab(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.cin(gnd),
	.combout(\Mux12~2_combout ),
	.cout());
defparam \Mux12~2 .lut_mask = 16'hFFDE;
defparam \Mux12~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux12~3 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datac(\Mux12~2_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.cin(gnd),
	.combout(\Mux12~3_combout ),
	.cout());
defparam \Mux12~3 .lut_mask = 16'hFFBE;
defparam \Mux12~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux12~4 (
	.dataa(\Mux12~1_combout ),
	.datab(\Mux12~3_combout ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ),
	.cin(gnd),
	.combout(\Mux12~4_combout ),
	.cout());
defparam \Mux12~4 .lut_mask = 16'hACFF;
defparam \Mux12~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux12~5 (
	.dataa(\Mux12~4_combout ),
	.datab(\Mux0~0_combout ),
	.datac(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux12~5_combout ),
	.cout());
defparam \Mux12~5 .lut_mask = 16'hFEFE;
defparam \Mux12~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux11~0 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datab(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
defparam \Mux11~0 .lut_mask = 16'hFFDE;
defparam \Mux11~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux11~1 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datac(\Mux11~0_combout ),
	.datad(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.cin(gnd),
	.combout(\Mux11~1_combout ),
	.cout());
defparam \Mux11~1 .lut_mask = 16'hFFBE;
defparam \Mux11~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux11~2 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datab(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.cin(gnd),
	.combout(\Mux11~2_combout ),
	.cout());
defparam \Mux11~2 .lut_mask = 16'hFFDE;
defparam \Mux11~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux11~3 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datac(\Mux11~2_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.cin(gnd),
	.combout(\Mux11~3_combout ),
	.cout());
defparam \Mux11~3 .lut_mask = 16'hFFBE;
defparam \Mux11~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux11~4 (
	.dataa(\Mux11~1_combout ),
	.datab(\Mux11~3_combout ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ),
	.cin(gnd),
	.combout(\Mux11~4_combout ),
	.cout());
defparam \Mux11~4 .lut_mask = 16'hACFF;
defparam \Mux11~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux11~5 (
	.dataa(\Mux11~4_combout ),
	.datab(\Mux0~0_combout ),
	.datac(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux11~5_combout ),
	.cout());
defparam \Mux11~5 .lut_mask = 16'hFEFE;
defparam \Mux11~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux10~0 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datab(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
defparam \Mux10~0 .lut_mask = 16'hFFDE;
defparam \Mux10~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux10~1 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datac(\Mux10~0_combout ),
	.datad(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.cin(gnd),
	.combout(\Mux10~1_combout ),
	.cout());
defparam \Mux10~1 .lut_mask = 16'hFFBE;
defparam \Mux10~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux10~2 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datab(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.cin(gnd),
	.combout(\Mux10~2_combout ),
	.cout());
defparam \Mux10~2 .lut_mask = 16'hFFDE;
defparam \Mux10~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux10~3 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datac(\Mux10~2_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.cin(gnd),
	.combout(\Mux10~3_combout ),
	.cout());
defparam \Mux10~3 .lut_mask = 16'hFFBE;
defparam \Mux10~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux10~4 (
	.dataa(\Mux10~1_combout ),
	.datab(\Mux10~3_combout ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ),
	.cin(gnd),
	.combout(\Mux10~4_combout ),
	.cout());
defparam \Mux10~4 .lut_mask = 16'hACFF;
defparam \Mux10~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux10~5 (
	.dataa(\Mux10~4_combout ),
	.datab(\Mux0~0_combout ),
	.datac(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux10~5_combout ),
	.cout());
defparam \Mux10~5 .lut_mask = 16'hFEFE;
defparam \Mux10~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux9~0 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datab(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
defparam \Mux9~0 .lut_mask = 16'hFFDE;
defparam \Mux9~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux9~1 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datac(\Mux9~0_combout ),
	.datad(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.cin(gnd),
	.combout(\Mux9~1_combout ),
	.cout());
defparam \Mux9~1 .lut_mask = 16'hFFBE;
defparam \Mux9~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux9~2 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datab(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.cin(gnd),
	.combout(\Mux9~2_combout ),
	.cout());
defparam \Mux9~2 .lut_mask = 16'hFFDE;
defparam \Mux9~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux9~3 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datac(\Mux9~2_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.cin(gnd),
	.combout(\Mux9~3_combout ),
	.cout());
defparam \Mux9~3 .lut_mask = 16'hFFBE;
defparam \Mux9~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux9~4 (
	.dataa(\Mux9~1_combout ),
	.datab(\Mux9~3_combout ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ),
	.cin(gnd),
	.combout(\Mux9~4_combout ),
	.cout());
defparam \Mux9~4 .lut_mask = 16'hACFF;
defparam \Mux9~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux9~5 (
	.dataa(\Mux9~4_combout ),
	.datab(\Mux0~0_combout ),
	.datac(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux9~5_combout ),
	.cout());
defparam \Mux9~5 .lut_mask = 16'hFEFE;
defparam \Mux9~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux8~0 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datab(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
defparam \Mux8~0 .lut_mask = 16'hFFDE;
defparam \Mux8~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux8~1 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datac(\Mux8~0_combout ),
	.datad(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.cin(gnd),
	.combout(\Mux8~1_combout ),
	.cout());
defparam \Mux8~1 .lut_mask = 16'hFFBE;
defparam \Mux8~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux8~2 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datab(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.cin(gnd),
	.combout(\Mux8~2_combout ),
	.cout());
defparam \Mux8~2 .lut_mask = 16'hFFDE;
defparam \Mux8~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux8~3 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datac(\Mux8~2_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.cin(gnd),
	.combout(\Mux8~3_combout ),
	.cout());
defparam \Mux8~3 .lut_mask = 16'hFFBE;
defparam \Mux8~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux8~4 (
	.dataa(\Mux8~1_combout ),
	.datab(\Mux8~3_combout ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ),
	.cin(gnd),
	.combout(\Mux8~4_combout ),
	.cout());
defparam \Mux8~4 .lut_mask = 16'hACFF;
defparam \Mux8~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux8~5 (
	.dataa(\Mux8~4_combout ),
	.datab(\Mux0~0_combout ),
	.datac(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux8~5_combout ),
	.cout());
defparam \Mux8~5 .lut_mask = 16'hFEFE;
defparam \Mux8~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux7~0 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datab(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
defparam \Mux7~0 .lut_mask = 16'hFFDE;
defparam \Mux7~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux7~1 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datac(\Mux7~0_combout ),
	.datad(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
defparam \Mux7~1 .lut_mask = 16'hFFBE;
defparam \Mux7~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux7~2 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datab(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.cin(gnd),
	.combout(\Mux7~2_combout ),
	.cout());
defparam \Mux7~2 .lut_mask = 16'hFFDE;
defparam \Mux7~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux7~3 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datac(\Mux7~2_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.cin(gnd),
	.combout(\Mux7~3_combout ),
	.cout());
defparam \Mux7~3 .lut_mask = 16'hFFBE;
defparam \Mux7~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux7~4 (
	.dataa(\Mux7~1_combout ),
	.datab(\Mux7~3_combout ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ),
	.cin(gnd),
	.combout(\Mux7~4_combout ),
	.cout());
defparam \Mux7~4 .lut_mask = 16'hACFF;
defparam \Mux7~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux7~5 (
	.dataa(\Mux7~4_combout ),
	.datab(\Mux0~0_combout ),
	.datac(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux7~5_combout ),
	.cout());
defparam \Mux7~5 .lut_mask = 16'hFEFE;
defparam \Mux7~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux6~0 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datab(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
defparam \Mux6~0 .lut_mask = 16'hFFDE;
defparam \Mux6~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux6~1 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datac(\Mux6~0_combout ),
	.datad(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
defparam \Mux6~1 .lut_mask = 16'hFFBE;
defparam \Mux6~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux6~2 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datab(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.cin(gnd),
	.combout(\Mux6~2_combout ),
	.cout());
defparam \Mux6~2 .lut_mask = 16'hFFDE;
defparam \Mux6~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux6~3 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datac(\Mux6~2_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.cin(gnd),
	.combout(\Mux6~3_combout ),
	.cout());
defparam \Mux6~3 .lut_mask = 16'hFFBE;
defparam \Mux6~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux6~4 (
	.dataa(\Mux6~1_combout ),
	.datab(\Mux6~3_combout ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ),
	.cin(gnd),
	.combout(\Mux6~4_combout ),
	.cout());
defparam \Mux6~4 .lut_mask = 16'hACFF;
defparam \Mux6~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux6~5 (
	.dataa(\Mux6~4_combout ),
	.datab(\Mux0~0_combout ),
	.datac(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux6~5_combout ),
	.cout());
defparam \Mux6~5 .lut_mask = 16'hFEFE;
defparam \Mux6~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux5~0 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datab(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
defparam \Mux5~0 .lut_mask = 16'hFFDE;
defparam \Mux5~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux5~1 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datac(\Mux5~0_combout ),
	.datad(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
defparam \Mux5~1 .lut_mask = 16'hFFBE;
defparam \Mux5~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux5~2 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datab(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.cin(gnd),
	.combout(\Mux5~2_combout ),
	.cout());
defparam \Mux5~2 .lut_mask = 16'hFFDE;
defparam \Mux5~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux5~3 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datac(\Mux5~2_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.cin(gnd),
	.combout(\Mux5~3_combout ),
	.cout());
defparam \Mux5~3 .lut_mask = 16'hFFBE;
defparam \Mux5~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux5~4 (
	.dataa(\Mux5~1_combout ),
	.datab(\Mux5~3_combout ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ),
	.cin(gnd),
	.combout(\Mux5~4_combout ),
	.cout());
defparam \Mux5~4 .lut_mask = 16'hACFF;
defparam \Mux5~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux5~5 (
	.dataa(\Mux5~4_combout ),
	.datab(\Mux0~0_combout ),
	.datac(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux5~5_combout ),
	.cout());
defparam \Mux5~5 .lut_mask = 16'hFEFE;
defparam \Mux5~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux4~0 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datab(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
defparam \Mux4~0 .lut_mask = 16'hFFDE;
defparam \Mux4~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux4~1 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datac(\Mux4~0_combout ),
	.datad(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
defparam \Mux4~1 .lut_mask = 16'hFFBE;
defparam \Mux4~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux4~2 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datab(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.cin(gnd),
	.combout(\Mux4~2_combout ),
	.cout());
defparam \Mux4~2 .lut_mask = 16'hFFDE;
defparam \Mux4~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux4~3 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datac(\Mux4~2_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.cin(gnd),
	.combout(\Mux4~3_combout ),
	.cout());
defparam \Mux4~3 .lut_mask = 16'hFFBE;
defparam \Mux4~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux4~4 (
	.dataa(\Mux4~1_combout ),
	.datab(\Mux4~3_combout ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ),
	.cin(gnd),
	.combout(\Mux4~4_combout ),
	.cout());
defparam \Mux4~4 .lut_mask = 16'hACFF;
defparam \Mux4~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux4~5 (
	.dataa(\Mux4~4_combout ),
	.datab(\Mux0~0_combout ),
	.datac(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux4~5_combout ),
	.cout());
defparam \Mux4~5 .lut_mask = 16'hFEFE;
defparam \Mux4~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux3~0 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datab(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'hFFDE;
defparam \Mux3~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux3~1 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datac(\Mux3~0_combout ),
	.datad(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
defparam \Mux3~1 .lut_mask = 16'hFFBE;
defparam \Mux3~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux3~2 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datab(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.cin(gnd),
	.combout(\Mux3~2_combout ),
	.cout());
defparam \Mux3~2 .lut_mask = 16'hFFDE;
defparam \Mux3~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux3~3 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datac(\Mux3~2_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.cin(gnd),
	.combout(\Mux3~3_combout ),
	.cout());
defparam \Mux3~3 .lut_mask = 16'hFFBE;
defparam \Mux3~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux3~4 (
	.dataa(\Mux3~1_combout ),
	.datab(\Mux3~3_combout ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ),
	.cin(gnd),
	.combout(\Mux3~4_combout ),
	.cout());
defparam \Mux3~4 .lut_mask = 16'hACFF;
defparam \Mux3~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux3~5 (
	.dataa(\Mux3~4_combout ),
	.datab(\Mux0~0_combout ),
	.datac(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux3~5_combout ),
	.cout());
defparam \Mux3~5 .lut_mask = 16'hFEFE;
defparam \Mux3~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux2~0 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datab(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hFFDE;
defparam \Mux2~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux2~1 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datac(\Mux2~0_combout ),
	.datad(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
defparam \Mux2~1 .lut_mask = 16'hFFBE;
defparam \Mux2~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux2~2 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datab(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.cin(gnd),
	.combout(\Mux2~2_combout ),
	.cout());
defparam \Mux2~2 .lut_mask = 16'hFFDE;
defparam \Mux2~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux2~3 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datac(\Mux2~2_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.cin(gnd),
	.combout(\Mux2~3_combout ),
	.cout());
defparam \Mux2~3 .lut_mask = 16'hFFBE;
defparam \Mux2~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux2~4 (
	.dataa(\Mux2~1_combout ),
	.datab(\Mux2~3_combout ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ),
	.cin(gnd),
	.combout(\Mux2~4_combout ),
	.cout());
defparam \Mux2~4 .lut_mask = 16'hACFF;
defparam \Mux2~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux2~5 (
	.dataa(\Mux2~4_combout ),
	.datab(\Mux0~0_combout ),
	.datac(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux2~5_combout ),
	.cout());
defparam \Mux2~5 .lut_mask = 16'hFEFE;
defparam \Mux2~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux1~0 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datab(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hFFDE;
defparam \Mux1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux1~1 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datac(\Mux1~0_combout ),
	.datad(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hFFBE;
defparam \Mux1~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux1~2 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datab(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
defparam \Mux1~2 .lut_mask = 16'hFFDE;
defparam \Mux1~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux1~3 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datac(\Mux1~2_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.cin(gnd),
	.combout(\Mux1~3_combout ),
	.cout());
defparam \Mux1~3 .lut_mask = 16'hFFBE;
defparam \Mux1~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux1~4 (
	.dataa(\Mux1~1_combout ),
	.datab(\Mux1~3_combout ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ),
	.cin(gnd),
	.combout(\Mux1~4_combout ),
	.cout());
defparam \Mux1~4 .lut_mask = 16'hACFF;
defparam \Mux1~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux1~5 (
	.dataa(\Mux1~4_combout ),
	.datab(\Mux0~0_combout ),
	.datac(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux1~5_combout ),
	.cout());
defparam \Mux1~5 .lut_mask = 16'hFEFE;
defparam \Mux1~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux0~1 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datab(\integrator[6].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datad(\integrator[4].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hFFDE;
defparam \Mux0~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux0~2 (
	.dataa(\integrator[5].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datac(\Mux0~1_combout ),
	.datad(\integrator[7].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
defparam \Mux0~2 .lut_mask = 16'hFFBE;
defparam \Mux0~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux0~3 (
	.dataa(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datab(\integrator[1].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[155]~8_combout ),
	.datad(\integrator[0].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
defparam \Mux0~3 .lut_mask = 16'hFFDE;
defparam \Mux0~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux0~4 (
	.dataa(\integrator[2].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.datab(\Mod2|auto_generated|divider|divider|StageOut[156]~9_combout ),
	.datac(\Mux0~3_combout ),
	.datad(\integrator[3].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.cin(gnd),
	.combout(\Mux0~4_combout ),
	.cout());
defparam \Mux0~4 .lut_mask = 16'hFFBE;
defparam \Mux0~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux0~5 (
	.dataa(\Mux0~2_combout ),
	.datab(\Mux0~4_combout ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[157]~10_combout ),
	.datad(\Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ),
	.cin(gnd),
	.combout(\Mux0~5_combout ),
	.cout());
defparam \Mux0~5 .lut_mask = 16'hACFF;
defparam \Mux0~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux0~6 (
	.dataa(\Mux0~5_combout ),
	.datab(\Mux0~0_combout ),
	.datac(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux0~6_combout ),
	.cout());
defparam \Mux0~6 .lut_mask = 16'hFEFE;
defparam \Mux0~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \ena_diff_s~1 (
	.dataa(reset_n),
	.datab(\ena_sample~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ena_diff_s~1_combout ),
	.cout());
defparam \ena_diff_s~1 .lut_mask = 16'hEEEE;
defparam \ena_diff_s~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \ena_sample~0 (
	.dataa(\sample_state[0]~q ),
	.datab(gnd),
	.datac(stall_reg),
	.datad(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[6]~q ),
	.cin(gnd),
	.combout(\ena_sample~0_combout ),
	.cout());
defparam \ena_sample~0 .lut_mask = 16'hAFFF;
defparam \ena_sample~0 .sum_lutc_input = "datac";

dffeas \fifo_rdreq[5] (
	.clk(clk),
	.d(\always5~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[5]~q ),
	.prn(vcc));
defparam \fifo_rdreq[5] .is_wysiwyg = "true";
defparam \fifo_rdreq[5] .power_up = "low";

dffeas \fifo_rdreq[6] (
	.clk(clk),
	.d(\always5~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[6]~q ),
	.prn(vcc));
defparam \fifo_rdreq[6] .is_wysiwyg = "true";
defparam \fifo_rdreq[6] .power_up = "low";

dffeas \fifo_rdreq[4] (
	.clk(clk),
	.d(\always5~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[4]~q ),
	.prn(vcc));
defparam \fifo_rdreq[4] .is_wysiwyg = "true";
defparam \fifo_rdreq[4] .power_up = "low";

dffeas \fifo_rdreq[7] (
	.clk(clk),
	.d(\always5~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[7]~q ),
	.prn(vcc));
defparam \fifo_rdreq[7] .is_wysiwyg = "true";
defparam \fifo_rdreq[7] .power_up = "low";

dffeas \fifo_rdreq[2] (
	.clk(clk),
	.d(\always5~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[2]~q ),
	.prn(vcc));
defparam \fifo_rdreq[2] .is_wysiwyg = "true";
defparam \fifo_rdreq[2] .power_up = "low";

dffeas \fifo_rdreq[1] (
	.clk(clk),
	.d(\always5~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[1]~q ),
	.prn(vcc));
defparam \fifo_rdreq[1] .is_wysiwyg = "true";
defparam \fifo_rdreq[1] .power_up = "low";

dffeas \fifo_rdreq[0] (
	.clk(clk),
	.d(\always5~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[0]~q ),
	.prn(vcc));
defparam \fifo_rdreq[0] .is_wysiwyg = "true";
defparam \fifo_rdreq[0] .power_up = "low";

dffeas \fifo_rdreq[3] (
	.clk(clk),
	.d(\always5~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[3]~q ),
	.prn(vcc));
defparam \fifo_rdreq[3] .is_wysiwyg = "true";
defparam \fifo_rdreq[3] .power_up = "low";

dffeas \fifo_rdreq[8] (
	.clk(clk),
	.d(\always5~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!stall_reg),
	.q(\fifo_rdreq[8]~q ),
	.prn(vcc));
defparam \fifo_rdreq[8] .is_wysiwyg = "true";
defparam \fifo_rdreq[8] .power_up = "low";

fiftyfivenm_lcell_comb \ena_sample~1 (
	.dataa(\ena_sample~q ),
	.datab(stall_reg),
	.datac(gnd),
	.datad(\sample_state[0]~q ),
	.cin(gnd),
	.combout(\ena_sample~1_combout ),
	.cout());
defparam \ena_sample~1 .lut_mask = 16'hEEFF;
defparam \ena_sample~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[10]~36 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[6]~q ),
	.datab(\Mod0|auto_generated|divider|divider|op_1~6_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[10]~36_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[10]~36 .lut_mask = 16'hEEEE;
defparam \Mod0|auto_generated|divider|divider|StageOut[10]~36 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[10]~37 (
	.dataa(\Mod0|auto_generated|divider|divider|op_1~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|op_1~6_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[10]~37_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[10]~37 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[10]~37 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[9]~38 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[5]~q ),
	.datab(\Mod0|auto_generated|divider|divider|op_1~6_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[9]~38_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[9]~38 .lut_mask = 16'hEEEE;
defparam \Mod0|auto_generated|divider|divider|StageOut[9]~38 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[9]~39 (
	.dataa(\Mod0|auto_generated|divider|divider|op_1~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|op_1~6_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[9]~39_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[9]~39 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[9]~39 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[8]~40 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[4]~q ),
	.datab(\Mod0|auto_generated|divider|divider|op_1~6_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[8]~40_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[8]~40 .lut_mask = 16'hEEEE;
defparam \Mod0|auto_generated|divider|divider|StageOut[8]~40 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[8]~41 (
	.dataa(\Mod0|auto_generated|divider|divider|op_1~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|op_1~6_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[8]~41_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[8]~41 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[8]~41 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[14]~42 (
	.dataa(\Mod0|auto_generated|divider|divider|op_2~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|op_2~8_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[14]~42_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[14]~42 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[14]~42 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[13]~43 (
	.dataa(\Mod0|auto_generated|divider|divider|op_2~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|op_2~8_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[13]~43_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[13]~43 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[13]~43 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[12]~44 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[3]~q ),
	.datab(\Mod0|auto_generated|divider|divider|op_2~8_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[12]~44_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[12]~44 .lut_mask = 16'hEEEE;
defparam \Mod0|auto_generated|divider|divider|StageOut[12]~44 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[12]~45 (
	.dataa(\Mod0|auto_generated|divider|divider|op_2~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|op_2~8_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[12]~45_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[12]~45 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[12]~45 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[18]~46 (
	.dataa(\Mod0|auto_generated|divider|divider|op_3~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|op_3~8_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[18]~46_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[18]~46 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[18]~46 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[17]~47 (
	.dataa(\Mod0|auto_generated|divider|divider|op_3~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|op_3~8_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[17]~47_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[17]~47 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[17]~47 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[16]~48 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[2]~q ),
	.datab(\Mod0|auto_generated|divider|divider|op_3~8_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[16]~48_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[16]~48 .lut_mask = 16'hEEEE;
defparam \Mod0|auto_generated|divider|divider|StageOut[16]~48 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[16]~49 (
	.dataa(\Mod0|auto_generated|divider|divider|op_3~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|op_3~8_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[16]~49_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[16]~49 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[16]~49 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[20]~50 (
	.dataa(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[1]~q ),
	.datab(\Mod0|auto_generated|divider|divider|op_4~8_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[20]~50_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[20]~50 .lut_mask = 16'hEEEE;
defparam \Mod0|auto_generated|divider|divider|StageOut[20]~50 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[20]~51 (
	.dataa(\Mod0|auto_generated|divider|divider|op_4~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|op_4~8_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[20]~51_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[20]~51 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[20]~51 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[21]~52 (
	.dataa(\Mod0|auto_generated|divider|divider|op_4~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|op_4~8_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[21]~52_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[21]~52 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[21]~52 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[22]~53 (
	.dataa(\Mod0|auto_generated|divider|divider|op_4~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mod0|auto_generated|divider|divider|op_4~8_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[22]~53_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[22]~53 .lut_mask = 16'hAAFF;
defparam \Mod0|auto_generated|divider|divider|StageOut[22]~53 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \ena_sample~2 (
	.dataa(\Mod0|auto_generated|divider|divider|op_5~0_combout ),
	.datab(\Mod0|auto_generated|divider|divider|op_5~2_combout ),
	.datac(\Mod0|auto_generated|divider|divider|op_5~4_combout ),
	.datad(\Mod0|auto_generated|divider|divider|op_5~8_combout ),
	.cin(gnd),
	.combout(\ena_sample~2_combout ),
	.cout());
defparam \ena_sample~2 .lut_mask = 16'h7FFF;
defparam \ena_sample~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \ena_sample~3 (
	.dataa(\Mod0|auto_generated|divider|divider|op_4~8_combout ),
	.datab(\Mod0|auto_generated|divider|divider|op_4~0_combout ),
	.datac(\Mod0|auto_generated|divider|divider|op_4~2_combout ),
	.datad(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[1]~q ),
	.cin(gnd),
	.combout(\ena_sample~3_combout ),
	.cout());
defparam \ena_sample~3 .lut_mask = 16'h27FF;
defparam \ena_sample~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \ena_sample~4 (
	.dataa(\Mod0|auto_generated|divider|divider|op_5~8_combout ),
	.datab(\ena_sample~3_combout ),
	.datac(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[0]~q ),
	.datad(\Mod0|auto_generated|divider|divider|StageOut[21]~59_combout ),
	.cin(gnd),
	.combout(\ena_sample~4_combout ),
	.cout());
defparam \ena_sample~4 .lut_mask = 16'hEFFF;
defparam \ena_sample~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \ena_sample~5 (
	.dataa(\ena_sample~1_combout ),
	.datab(\ena_sample~0_combout ),
	.datac(\ena_sample~2_combout ),
	.datad(\ena_sample~4_combout ),
	.cin(gnd),
	.combout(\ena_sample~5_combout ),
	.cout());
defparam \ena_sample~5 .lut_mask = 16'hFFFE;
defparam \ena_sample~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \sample_state~0 (
	.dataa(\latency_cnt[2]~q ),
	.datab(\latency_cnt[1]~q ),
	.datac(\latency_cnt[3]~q ),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\sample_state~0_combout ),
	.cout());
defparam \sample_state~0 .lut_mask = 16'hFEFF;
defparam \sample_state~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \sample_state~1 (
	.dataa(\sample_state[0]~q ),
	.datab(\sample_state~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sample_state~1_combout ),
	.cout());
defparam \sample_state~1 .lut_mask = 16'hEEEE;
defparam \sample_state~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod1|auto_generated|divider|divider|StageOut[12]~0 (
	.dataa(\int_channel_cnt_inst|count[0]~q ),
	.datab(\Mod1|auto_generated|divider|divider|op_2~0_combout ),
	.datac(gnd),
	.datad(\Mod1|auto_generated|divider|divider|op_2~8_combout ),
	.cin(gnd),
	.combout(\Mod1|auto_generated|divider|divider|StageOut[12]~0_combout ),
	.cout());
defparam \Mod1|auto_generated|divider|divider|StageOut[12]~0 .lut_mask = 16'hAACC;
defparam \Mod1|auto_generated|divider|divider|StageOut[12]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod1|auto_generated|divider|divider|StageOut[14]~1 (
	.dataa(\int_channel_cnt_inst|count[2]~q ),
	.datab(\Mod1|auto_generated|divider|divider|op_2~4_combout ),
	.datac(gnd),
	.datad(\Mod1|auto_generated|divider|divider|op_2~8_combout ),
	.cin(gnd),
	.combout(\Mod1|auto_generated|divider|divider|StageOut[14]~1_combout ),
	.cout());
defparam \Mod1|auto_generated|divider|divider|StageOut[14]~1 .lut_mask = 16'hAACC;
defparam \Mod1|auto_generated|divider|divider|StageOut[14]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \always5~0 (
	.dataa(\ena_sample~q ),
	.datab(\Mod1|auto_generated|divider|divider|op_2~8_combout ),
	.datac(\Mod1|auto_generated|divider|divider|op_2~6_combout ),
	.datad(\int_channel_cnt_inst|count[3]~q ),
	.cin(gnd),
	.combout(\always5~0_combout ),
	.cout());
defparam \always5~0 .lut_mask = 16'h8BFF;
defparam \always5~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod1|auto_generated|divider|divider|StageOut[13]~2 (
	.dataa(\int_channel_cnt_inst|count[1]~q ),
	.datab(\Mod1|auto_generated|divider|divider|op_2~2_combout ),
	.datac(gnd),
	.datad(\Mod1|auto_generated|divider|divider|op_2~8_combout ),
	.cin(gnd),
	.combout(\Mod1|auto_generated|divider|divider|StageOut[13]~2_combout ),
	.cout());
defparam \Mod1|auto_generated|divider|divider|StageOut[13]~2 .lut_mask = 16'hAACC;
defparam \Mod1|auto_generated|divider|divider|StageOut[13]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \always5~1 (
	.dataa(\Mod1|auto_generated|divider|divider|StageOut[12]~0_combout ),
	.datab(\Mod1|auto_generated|divider|divider|StageOut[14]~1_combout ),
	.datac(\always5~0_combout ),
	.datad(\Mod1|auto_generated|divider|divider|StageOut[13]~2_combout ),
	.cin(gnd),
	.combout(\always5~1_combout ),
	.cout());
defparam \always5~1 .lut_mask = 16'hFEFF;
defparam \always5~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \always5~2 (
	.dataa(\Mod1|auto_generated|divider|divider|StageOut[13]~2_combout ),
	.datab(\Mod1|auto_generated|divider|divider|StageOut[14]~1_combout ),
	.datac(\always5~0_combout ),
	.datad(\Mod1|auto_generated|divider|divider|StageOut[12]~0_combout ),
	.cin(gnd),
	.combout(\always5~2_combout ),
	.cout());
defparam \always5~2 .lut_mask = 16'hFEFF;
defparam \always5~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \always5~3 (
	.dataa(\Mod1|auto_generated|divider|divider|StageOut[14]~1_combout ),
	.datab(\always5~0_combout ),
	.datac(\Mod1|auto_generated|divider|divider|StageOut[13]~2_combout ),
	.datad(\Mod1|auto_generated|divider|divider|StageOut[12]~0_combout ),
	.cin(gnd),
	.combout(\always5~3_combout ),
	.cout());
defparam \always5~3 .lut_mask = 16'hEFFF;
defparam \always5~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \always5~4 (
	.dataa(\Mod1|auto_generated|divider|divider|StageOut[13]~2_combout ),
	.datab(\Mod1|auto_generated|divider|divider|StageOut[12]~0_combout ),
	.datac(\Mod1|auto_generated|divider|divider|StageOut[14]~1_combout ),
	.datad(\always5~0_combout ),
	.cin(gnd),
	.combout(\always5~4_combout ),
	.cout());
defparam \always5~4 .lut_mask = 16'hFFFE;
defparam \always5~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \always5~5 (
	.dataa(\Mod1|auto_generated|divider|divider|StageOut[13]~2_combout ),
	.datab(\always5~0_combout ),
	.datac(\Mod1|auto_generated|divider|divider|StageOut[12]~0_combout ),
	.datad(\Mod1|auto_generated|divider|divider|StageOut[14]~1_combout ),
	.cin(gnd),
	.combout(\always5~5_combout ),
	.cout());
defparam \always5~5 .lut_mask = 16'hEFFF;
defparam \always5~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \always5~6 (
	.dataa(\Mod1|auto_generated|divider|divider|StageOut[12]~0_combout ),
	.datab(\always5~0_combout ),
	.datac(\Mod1|auto_generated|divider|divider|StageOut[13]~2_combout ),
	.datad(\Mod1|auto_generated|divider|divider|StageOut[14]~1_combout ),
	.cin(gnd),
	.combout(\always5~6_combout ),
	.cout());
defparam \always5~6 .lut_mask = 16'hEFFF;
defparam \always5~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \always5~7 (
	.dataa(\always5~0_combout ),
	.datab(\Mod1|auto_generated|divider|divider|StageOut[13]~2_combout ),
	.datac(\Mod1|auto_generated|divider|divider|StageOut[12]~0_combout ),
	.datad(\Mod1|auto_generated|divider|divider|StageOut[14]~1_combout ),
	.cin(gnd),
	.combout(\always5~7_combout ),
	.cout());
defparam \always5~7 .lut_mask = 16'hBFFF;
defparam \always5~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \always5~8 (
	.dataa(\Mod1|auto_generated|divider|divider|StageOut[13]~2_combout ),
	.datab(\Mod1|auto_generated|divider|divider|StageOut[12]~0_combout ),
	.datac(\always5~0_combout ),
	.datad(\Mod1|auto_generated|divider|divider|StageOut[14]~1_combout ),
	.cin(gnd),
	.combout(\always5~8_combout ),
	.cout());
defparam \always5~8 .lut_mask = 16'hFEFF;
defparam \always5~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \always5~9 (
	.dataa(\ena_sample~q ),
	.datab(\int_channel_cnt_inst|count[3]~q ),
	.datac(\Mod1|auto_generated|divider|divider|op_2~6_combout ),
	.datad(\Mod1|auto_generated|divider|divider|op_2~8_combout ),
	.cin(gnd),
	.combout(\always5~9_combout ),
	.cout());
defparam \always5~9 .lut_mask = 16'hFAFC;
defparam \always5~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \always5~10 (
	.dataa(\always5~9_combout ),
	.datab(\Mod1|auto_generated|divider|divider|StageOut[13]~2_combout ),
	.datac(\Mod1|auto_generated|divider|divider|StageOut[12]~0_combout ),
	.datad(\Mod1|auto_generated|divider|divider|StageOut[14]~1_combout ),
	.cin(gnd),
	.combout(\always5~10_combout ),
	.cout());
defparam \always5~10 .lut_mask = 16'hBFFF;
defparam \always5~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux17~7 (
	.dataa(\Mux0~0_combout ),
	.datab(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ),
	.datad(\Mux17~6_combout ),
	.cin(gnd),
	.combout(\Mux17~7_combout ),
	.cout());
defparam \Mux17~7 .lut_mask = 16'hFFEF;
defparam \Mux17~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux16~7 (
	.dataa(\Mux0~0_combout ),
	.datab(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ),
	.datad(\Mux16~6_combout ),
	.cin(gnd),
	.combout(\Mux16~7_combout ),
	.cout());
defparam \Mux16~7 .lut_mask = 16'hFFEF;
defparam \Mux16~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux15~7 (
	.dataa(\Mux0~0_combout ),
	.datab(\integrator[8].fifo_regulator|buffer_FIFO|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.datac(\Mod2|auto_generated|divider|divider|StageOut[158]~11_combout ),
	.datad(\Mux15~6_combout ),
	.cin(gnd),
	.combout(\Mux15~7_combout ),
	.cout());
defparam \Mux15~7 .lut_mask = 16'hFFEF;
defparam \Mux15~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[18]~54 (
	.dataa(\Mod0|auto_generated|divider|divider|op_2~2_combout ),
	.datab(\Mod0|auto_generated|divider|divider|op_2~8_combout ),
	.datac(\Mod0|auto_generated|divider|divider|op_3~8_combout ),
	.datad(\Mod0|auto_generated|divider|divider|StageOut[13]~57_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[18]~54_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[18]~54 .lut_mask = 16'hFFFB;
defparam \Mod0|auto_generated|divider|divider|StageOut[18]~54 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[22]~55 (
	.dataa(\Mod0|auto_generated|divider|divider|op_3~2_combout ),
	.datab(\Mod0|auto_generated|divider|divider|op_3~8_combout ),
	.datac(\Mod0|auto_generated|divider|divider|op_4~8_combout ),
	.datad(\Mod0|auto_generated|divider|divider|StageOut[17]~58_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[22]~55_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[22]~55 .lut_mask = 16'hFFFB;
defparam \Mod0|auto_generated|divider|divider|StageOut[22]~55 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[14]~56 (
	.dataa(\Mod0|auto_generated|divider|divider|op_1~2_combout ),
	.datab(\Mod0|auto_generated|divider|divider|op_1~6_combout ),
	.datac(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[5]~q ),
	.datad(\Mod0|auto_generated|divider|divider|op_2~8_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[14]~56_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[14]~56 .lut_mask = 16'hFFB8;
defparam \Mod0|auto_generated|divider|divider|StageOut[14]~56 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[13]~57 (
	.dataa(\Mod0|auto_generated|divider|divider|op_1~0_combout ),
	.datab(\Mod0|auto_generated|divider|divider|op_1~6_combout ),
	.datac(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[4]~q ),
	.datad(\Mod0|auto_generated|divider|divider|op_2~8_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[13]~57_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[13]~57 .lut_mask = 16'hFFB8;
defparam \Mod0|auto_generated|divider|divider|StageOut[13]~57 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[17]~58 (
	.dataa(\Mod0|auto_generated|divider|divider|op_2~0_combout ),
	.datab(\Mod0|auto_generated|divider|divider|op_2~8_combout ),
	.datac(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[3]~q ),
	.datad(\Mod0|auto_generated|divider|divider|op_3~8_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[17]~58_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[17]~58 .lut_mask = 16'hFFB8;
defparam \Mod0|auto_generated|divider|divider|StageOut[17]~58 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mod0|auto_generated|divider|divider|StageOut[21]~59 (
	.dataa(\Mod0|auto_generated|divider|divider|op_3~0_combout ),
	.datab(\Mod0|auto_generated|divider|divider|op_3~8_combout ),
	.datac(\integrator[0].j0.vrc_en_0.first_dsample|counter_fs_inst|count[2]~q ),
	.datad(\Mod0|auto_generated|divider|divider|op_4~8_combout ),
	.cin(gnd),
	.combout(\Mod0|auto_generated|divider|divider|StageOut[21]~59_combout ),
	.cout());
defparam \Mod0|auto_generated|divider|divider|StageOut[21]~59 .lut_mask = 16'hFFB8;
defparam \Mod0|auto_generated|divider|divider|StageOut[21]~59 .sum_lutc_input = "datac";

dffeas \state[0] (
	.clk(clk),
	.d(\state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(state_0),
	.prn(vcc));
defparam \state[0] .is_wysiwyg = "true";
defparam \state[0] .power_up = "low";

dffeas \channel_out_int[3] (
	.clk(clk),
	.d(\channel_out_int~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\channel_out_int[1]~2_combout ),
	.q(channel_out_int_3),
	.prn(vcc));
defparam \channel_out_int[3] .is_wysiwyg = "true";
defparam \channel_out_int[3] .power_up = "low";

dffeas \channel_out_int[0] (
	.clk(clk),
	.d(\channel_out_int~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\channel_out_int[1]~2_combout ),
	.q(channel_out_int_0),
	.prn(vcc));
defparam \channel_out_int[0] .is_wysiwyg = "true";
defparam \channel_out_int[0] .power_up = "low";

dffeas \channel_out_int[1] (
	.clk(clk),
	.d(\channel_out_int~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\channel_out_int[1]~2_combout ),
	.q(channel_out_int_1),
	.prn(vcc));
defparam \channel_out_int[1] .is_wysiwyg = "true";
defparam \channel_out_int[1] .power_up = "low";

dffeas \channel_out_int[2] (
	.clk(clk),
	.d(\channel_out_int~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\channel_out_int[1]~2_combout ),
	.q(channel_out_int_2),
	.prn(vcc));
defparam \channel_out_int[2] .is_wysiwyg = "true";
defparam \channel_out_int[2] .power_up = "low";

fiftyfivenm_lcell_comb \latency_cnt[3]~0 (
	.dataa(reset_n),
	.datab(stall_reg),
	.datac(\state~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\latency_cnt[3]~0_combout ),
	.cout());
defparam \latency_cnt[3]~0 .lut_mask = 16'hFEFE;
defparam \latency_cnt[3]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \latency_cnt[0]~4 (
	.dataa(stall_reg),
	.datab(\latency_cnt[0]~q ),
	.datac(\state~0_combout ),
	.datad(reset_n),
	.cin(gnd),
	.combout(\latency_cnt[0]~4_combout ),
	.cout());
defparam \latency_cnt[0]~4 .lut_mask = 16'h6FFF;
defparam \latency_cnt[0]~4 .sum_lutc_input = "datac";

dffeas \latency_cnt[0] (
	.clk(clk),
	.d(\latency_cnt[0]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\latency_cnt[0]~q ),
	.prn(vcc));
defparam \latency_cnt[0] .is_wysiwyg = "true";
defparam \latency_cnt[0] .power_up = "low";

fiftyfivenm_lcell_comb \latency_cnt[1]~3 (
	.dataa(\latency_cnt[1]~q ),
	.datab(\latency_cnt[3]~0_combout ),
	.datac(reset_n),
	.datad(\latency_cnt[0]~q ),
	.cin(gnd),
	.combout(\latency_cnt[1]~3_combout ),
	.cout());
defparam \latency_cnt[1]~3 .lut_mask = 16'hF9F6;
defparam \latency_cnt[1]~3 .sum_lutc_input = "datac";

dffeas \latency_cnt[1] (
	.clk(clk),
	.d(\latency_cnt[1]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\latency_cnt[1]~q ),
	.prn(vcc));
defparam \latency_cnt[1] .is_wysiwyg = "true";
defparam \latency_cnt[1] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~1 (
	.dataa(gnd),
	.datab(\latency_cnt[2]~q ),
	.datac(\latency_cnt[1]~q ),
	.datad(\latency_cnt[0]~q ),
	.cin(gnd),
	.combout(\Add3~1_combout ),
	.cout());
defparam \Add3~1 .lut_mask = 16'hC33C;
defparam \Add3~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \latency_cnt[2]~2 (
	.dataa(\latency_cnt[2]~q ),
	.datab(reset_n),
	.datac(\Add3~1_combout ),
	.datad(\latency_cnt[3]~0_combout ),
	.cin(gnd),
	.combout(\latency_cnt[2]~2_combout ),
	.cout());
defparam \latency_cnt[2]~2 .lut_mask = 16'hFAFC;
defparam \latency_cnt[2]~2 .sum_lutc_input = "datac";

dffeas \latency_cnt[2] (
	.clk(clk),
	.d(\latency_cnt[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\latency_cnt[2]~q ),
	.prn(vcc));
defparam \latency_cnt[2] .is_wysiwyg = "true";
defparam \latency_cnt[2] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~0 (
	.dataa(\latency_cnt[3]~q ),
	.datab(\latency_cnt[2]~q ),
	.datac(\latency_cnt[1]~q ),
	.datad(\latency_cnt[0]~q ),
	.cin(gnd),
	.combout(\Add3~0_combout ),
	.cout());
defparam \Add3~0 .lut_mask = 16'h6996;
defparam \Add3~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \latency_cnt[3]~1 (
	.dataa(\latency_cnt[3]~q ),
	.datab(reset_n),
	.datac(\Add3~0_combout ),
	.datad(\latency_cnt[3]~0_combout ),
	.cin(gnd),
	.combout(\latency_cnt[3]~1_combout ),
	.cout());
defparam \latency_cnt[3]~1 .lut_mask = 16'hFAFC;
defparam \latency_cnt[3]~1 .sum_lutc_input = "datac";

dffeas \latency_cnt[3] (
	.clk(clk),
	.d(\latency_cnt[3]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\latency_cnt[3]~q ),
	.prn(vcc));
defparam \latency_cnt[3] .is_wysiwyg = "true";
defparam \latency_cnt[3] .power_up = "low";

fiftyfivenm_lcell_comb \state~0 (
	.dataa(\latency_cnt[3]~q ),
	.datab(\latency_cnt[2]~q ),
	.datac(\latency_cnt[1]~q ),
	.datad(\latency_cnt[0]~q ),
	.cin(gnd),
	.combout(\state~0_combout ),
	.cout());
defparam \state~0 .lut_mask = 16'hBFFF;
defparam \state~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~1 (
	.dataa(state_0),
	.datab(\state~0_combout ),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\state~1_combout ),
	.cout());
defparam \state~1 .lut_mask = 16'hEEFF;
defparam \state~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~0 (
	.dataa(channel_out_int_3),
	.datab(channel_out_int_0),
	.datac(channel_out_int_1),
	.datad(channel_out_int_2),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
defparam \Add0~0 .lut_mask = 16'h6996;
defparam \Add0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \channel_out_int[1]~0 (
	.dataa(channel_out_int_0),
	.datab(channel_out_int_1),
	.datac(channel_out_int_2),
	.datad(channel_out_int_3),
	.cin(gnd),
	.combout(\channel_out_int[1]~0_combout ),
	.cout());
defparam \channel_out_int[1]~0 .lut_mask = 16'hFEFF;
defparam \channel_out_int[1]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \channel_out_int~1 (
	.dataa(reset_n),
	.datab(\Add0~0_combout ),
	.datac(\channel_out_int[1]~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\channel_out_int~1_combout ),
	.cout());
defparam \channel_out_int~1 .lut_mask = 16'hFEFE;
defparam \channel_out_int~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \channel_out_int[1]~2 (
	.dataa(reset_n),
	.datab(stall_reg),
	.datac(dout_valid),
	.datad(state_0),
	.cin(gnd),
	.combout(\channel_out_int[1]~2_combout ),
	.cout());
defparam \channel_out_int[1]~2 .lut_mask = 16'hFFF7;
defparam \channel_out_int[1]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \channel_out_int~3 (
	.dataa(channel_out_int_0),
	.datab(gnd),
	.datac(reset_n),
	.datad(\channel_out_int[1]~0_combout ),
	.cin(gnd),
	.combout(\channel_out_int~3_combout ),
	.cout());
defparam \channel_out_int~3 .lut_mask = 16'hFFF5;
defparam \channel_out_int~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \channel_out_int~4 (
	.dataa(reset_n),
	.datab(\channel_out_int[1]~0_combout ),
	.datac(channel_out_int_0),
	.datad(channel_out_int_1),
	.cin(gnd),
	.combout(\channel_out_int~4_combout ),
	.cout());
defparam \channel_out_int~4 .lut_mask = 16'hEFFE;
defparam \channel_out_int~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(channel_out_int_2),
	.datac(channel_out_int_0),
	.datad(channel_out_int_1),
	.cin(gnd),
	.combout(\Add0~1_combout ),
	.cout());
defparam \Add0~1 .lut_mask = 16'hC33C;
defparam \Add0~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \channel_out_int~5 (
	.dataa(reset_n),
	.datab(\channel_out_int[1]~0_combout ),
	.datac(\Add0~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\channel_out_int~5_combout ),
	.cout());
defparam \channel_out_int~5 .lut_mask = 16'hFEFE;
defparam \channel_out_int~5 .sum_lutc_input = "datac";

endmodule

module cic_auk_dspip_channel_buffer (
	q,
	count_1,
	count_2,
	count_3,
	count_4,
	count_0,
	count_5,
	data,
	stall_reg,
	ena_sample,
	valid_wreq,
	fifo_rdreq_0,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	count_1;
input 	count_2;
input 	count_3;
input 	count_4;
input 	count_0;
input 	count_5;
input 	[18:0] data;
input 	stall_reg;
input 	ena_sample;
output 	valid_wreq;
input 	fifo_rdreq_0;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_1 buffer_FIFO(
	.q({q_unconnected_wire_22,q_unconnected_wire_21,q_unconnected_wire_20,q_unconnected_wire_19,q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.count_1(count_1),
	.count_2(count_2),
	.count_3(count_3),
	.count_4(count_4),
	.count_0(count_0),
	.count_5(count_5),
	.data({gnd,gnd,gnd,gnd,data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.ena_sample(ena_sample),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_0(fifo_rdreq_0),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module cic_scfifo_1 (
	q,
	count_1,
	count_2,
	count_3,
	count_4,
	count_0,
	count_5,
	data,
	stall_reg,
	ena_sample,
	valid_wreq,
	fifo_rdreq_0,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[22:0] q;
input 	count_1;
input 	count_2;
input 	count_3;
input 	count_4;
input 	count_0;
input 	count_5;
input 	[22:0] data;
input 	stall_reg;
input 	ena_sample;
output 	valid_wreq;
input 	fifo_rdreq_0;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_1351 auto_generated(
	.q({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.count_1(count_1),
	.count_2(count_2),
	.count_3(count_3),
	.count_4(count_4),
	.count_0(count_0),
	.count_5(count_5),
	.data({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.ena_sample(ena_sample),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_0(fifo_rdreq_0),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module cic_scfifo_1351 (
	q,
	count_1,
	count_2,
	count_3,
	count_4,
	count_0,
	count_5,
	data,
	stall_reg,
	ena_sample,
	valid_wreq,
	fifo_rdreq_0,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	count_1;
input 	count_2;
input 	count_3;
input 	count_4;
input 	count_0;
input 	count_5;
input 	[18:0] data;
input 	stall_reg;
input 	ena_sample;
output 	valid_wreq;
input 	fifo_rdreq_0;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_a_dpfifo_c0u dpfifo(
	.q({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.count_1(count_1),
	.count_2(count_2),
	.count_3(count_3),
	.count_4(count_4),
	.count_0(count_0),
	.count_5(count_5),
	.data({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.ena_sample(ena_sample),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_0(fifo_rdreq_0),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module cic_a_dpfifo_c0u (
	q,
	count_1,
	count_2,
	count_3,
	count_4,
	count_0,
	count_5,
	data,
	stall_reg,
	ena_sample,
	valid_wreq,
	fifo_rdreq_0,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	count_1;
input 	count_2;
input 	count_3;
input 	count_4;
input 	count_0;
input 	count_5;
input 	[18:0] data;
input 	stall_reg;
input 	ena_sample;
output 	valid_wreq;
input 	fifo_rdreq_0;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \valid_wreq~2_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \empty_dff~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \valid_wreq~0_combout ;


cic_cntr_jka wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_cntr_vk6 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~2_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_cntr_ika rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_altsyncram_dlg1 FIFOram(
	.q_b({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data_a({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~2_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock0(clock),
	.clock1(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

fiftyfivenm_lcell_comb \valid_wreq~2 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~2_combout ),
	.cout());
defparam \valid_wreq~2 .lut_mask = 16'hAAFF;
defparam \valid_wreq~2 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

fiftyfivenm_lcell_comb \valid_rreq~0 (
	.dataa(fifo_rdreq_0),
	.datab(\empty_dff~q ),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(\usedw_counter|counter_reg_bit[3]~q ),
	.datac(\usedw_counter|counter_reg_bit[2]~q ),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hFEFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \_~1 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~0_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFEFF;
defparam \_~1 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

fiftyfivenm_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~2_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(\usedw_counter|counter_reg_bit[0]~q ),
	.datac(\usedw_counter|counter_reg_bit[3]~q ),
	.datad(\usedw_counter|counter_reg_bit[2]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~2 (
	.dataa(\usedw_will_be_1~1_combout ),
	.datab(\valid_wreq~2_combout ),
	.datac(\valid_rreq~0_combout ),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hEFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~2_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~1 (
	.dataa(fifo_rdreq_0),
	.datab(\empty_dff~q ),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hEEEE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \valid_wreq~1 (
	.dataa(ena_sample),
	.datab(\valid_wreq~0_combout ),
	.datac(count_0),
	.datad(count_5),
	.cin(gnd),
	.combout(valid_wreq),
	.cout());
defparam \valid_wreq~1 .lut_mask = 16'hEFFF;
defparam \valid_wreq~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \valid_wreq~0 (
	.dataa(count_1),
	.datab(count_2),
	.datac(count_3),
	.datad(count_4),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'h7FFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

endmodule

module cic_altsyncram_dlg1 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q_b;
input 	[18:0] data_a;
input 	[3:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[3:0] address_b;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

fiftyfivenm_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk1_output_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 19;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 19;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk1_output_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 19;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 19;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk1_output_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 19;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 19;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk1_output_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 19;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 19;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk1_output_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 19;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 19;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 19;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 19;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 19;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 19;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 19;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 19;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 19;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 19;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 19;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 19;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 19;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 19;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 19;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 19;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 19;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 19;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 19;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 19;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 19;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 19;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 19;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 19;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 4;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 15;
defparam ram_block1a16.port_a_logical_ram_depth = 16;
defparam ram_block1a16.port_a_logical_ram_width = 19;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 4;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 15;
defparam ram_block1a16.port_b_logical_ram_depth = 16;
defparam ram_block1a16.port_b_logical_ram_width = 19;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 4;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 15;
defparam ram_block1a17.port_a_logical_ram_depth = 16;
defparam ram_block1a17.port_a_logical_ram_width = 19;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 4;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 15;
defparam ram_block1a17.port_b_logical_ram_depth = 16;
defparam ram_block1a17.port_b_logical_ram_width = 19;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[0].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 4;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 15;
defparam ram_block1a18.port_a_logical_ram_depth = 16;
defparam ram_block1a18.port_a_logical_ram_width = 19;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 4;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 15;
defparam ram_block1a18.port_b_logical_ram_depth = 16;
defparam ram_block1a18.port_b_logical_ram_width = 19;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

endmodule

module cic_cntr_ika (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout());
defparam counter_comb_bita2.lut_mask = 16'h5A5A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

endmodule

module cic_cntr_jka (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module cic_cntr_vk6 (
	full_dff,
	counter_reg_bit_1,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_0,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_1;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_0;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_channel_buffer_1 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_1,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_1;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_2 buffer_FIFO(
	.q({q_unconnected_wire_22,q_unconnected_wire_21,q_unconnected_wire_20,q_unconnected_wire_19,q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({gnd,gnd,gnd,gnd,data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_1(fifo_rdreq_1),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module cic_scfifo_2 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_1,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[22:0] q;
input 	[22:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_1;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_1351_1 auto_generated(
	.q({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_1(fifo_rdreq_1),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module cic_scfifo_1351_1 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_1,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_1;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_a_dpfifo_c0u_1 dpfifo(
	.q({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_1(fifo_rdreq_1),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module cic_a_dpfifo_c0u_1 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_1,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_1;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \empty_dff~2_combout ;


cic_cntr_jka_1 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_cntr_vk6_1 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_cntr_ika_1 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_altsyncram_dlg1_1 FIFOram(
	.q_b({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data_a({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock0(clock),
	.clock1(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

fiftyfivenm_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

fiftyfivenm_lcell_comb \valid_rreq~0 (
	.dataa(fifo_rdreq_1),
	.datab(\empty_dff~q ),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(\usedw_counter|counter_reg_bit[3]~q ),
	.datac(\usedw_counter|counter_reg_bit[2]~q ),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hFEFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \_~1 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~0_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFEFF;
defparam \_~1 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

fiftyfivenm_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(\usedw_counter|counter_reg_bit[0]~q ),
	.datac(\usedw_counter|counter_reg_bit[3]~q ),
	.datad(\usedw_counter|counter_reg_bit[2]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~2 (
	.dataa(stall_reg),
	.datab(fifo_rdreq_1),
	.datac(\empty_dff~q ),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFFFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~1 (
	.dataa(fifo_rdreq_1),
	.datab(\empty_dff~q ),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

endmodule

module cic_altsyncram_dlg1_1 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q_b;
input 	[18:0] data_a;
input 	[3:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[3:0] address_b;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

fiftyfivenm_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk1_output_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 19;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 19;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk1_output_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 19;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 19;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk1_output_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 19;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 19;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk1_output_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 19;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 19;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk1_output_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 19;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 19;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 19;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 19;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 19;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 19;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 19;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 19;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 19;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 19;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 19;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 19;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 19;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 19;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 19;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 19;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 19;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 19;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 19;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 19;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 19;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 19;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 19;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 19;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 4;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 15;
defparam ram_block1a16.port_a_logical_ram_depth = 16;
defparam ram_block1a16.port_a_logical_ram_width = 19;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 4;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 15;
defparam ram_block1a16.port_b_logical_ram_depth = 16;
defparam ram_block1a16.port_b_logical_ram_width = 19;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 4;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 15;
defparam ram_block1a17.port_a_logical_ram_depth = 16;
defparam ram_block1a17.port_a_logical_ram_width = 19;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 4;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 15;
defparam ram_block1a17.port_b_logical_ram_depth = 16;
defparam ram_block1a17.port_b_logical_ram_width = 19;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[1].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 4;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 15;
defparam ram_block1a18.port_a_logical_ram_depth = 16;
defparam ram_block1a18.port_a_logical_ram_width = 19;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 4;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 15;
defparam ram_block1a18.port_b_logical_ram_depth = 16;
defparam ram_block1a18.port_b_logical_ram_width = 19;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

endmodule

module cic_cntr_ika_1 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout());
defparam counter_comb_bita2.lut_mask = 16'h5A5A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

endmodule

module cic_cntr_jka_1 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module cic_cntr_vk6_1 (
	full_dff,
	counter_reg_bit_1,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_0,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_1;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_0;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_channel_buffer_2 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_2,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_2;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_3 buffer_FIFO(
	.q({q_unconnected_wire_22,q_unconnected_wire_21,q_unconnected_wire_20,q_unconnected_wire_19,q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({gnd,gnd,gnd,gnd,data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_2(fifo_rdreq_2),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module cic_scfifo_3 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_2,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[22:0] q;
input 	[22:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_2;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_1351_2 auto_generated(
	.q({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_2(fifo_rdreq_2),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module cic_scfifo_1351_2 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_2,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_2;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_a_dpfifo_c0u_2 dpfifo(
	.q({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_2(fifo_rdreq_2),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module cic_a_dpfifo_c0u_2 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_2,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_2;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \empty_dff~2_combout ;
wire \usedw_will_be_1~3_combout ;


cic_cntr_jka_2 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_cntr_vk6_2 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_cntr_ika_2 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_altsyncram_dlg1_2 FIFOram(
	.q_b({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data_a({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock0(clock),
	.clock1(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

fiftyfivenm_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

fiftyfivenm_lcell_comb \valid_rreq~0 (
	.dataa(fifo_rdreq_2),
	.datab(\empty_dff~q ),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(\usedw_counter|counter_reg_bit[3]~q ),
	.datac(\usedw_counter|counter_reg_bit[2]~q ),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hFEFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \_~1 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~0_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFEFF;
defparam \_~1 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

fiftyfivenm_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(\usedw_counter|counter_reg_bit[0]~q ),
	.datac(\usedw_counter|counter_reg_bit[3]~q ),
	.datad(\usedw_counter|counter_reg_bit[2]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~2 (
	.dataa(\usedw_will_be_1~1_combout ),
	.datab(\valid_wreq~0_combout ),
	.datac(\valid_rreq~0_combout ),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hEFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~1 (
	.dataa(fifo_rdreq_2),
	.datab(\empty_dff~q ),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hEEEE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

endmodule

module cic_altsyncram_dlg1_2 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q_b;
input 	[18:0] data_a;
input 	[3:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[3:0] address_b;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

fiftyfivenm_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk1_output_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 19;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 19;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk1_output_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 19;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 19;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk1_output_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 19;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 19;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk1_output_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 19;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 19;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk1_output_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 19;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 19;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 19;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 19;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 19;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 19;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 19;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 19;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 19;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 19;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 19;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 19;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 19;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 19;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 19;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 19;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 19;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 19;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 19;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 19;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 19;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 19;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 19;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 19;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 4;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 15;
defparam ram_block1a16.port_a_logical_ram_depth = 16;
defparam ram_block1a16.port_a_logical_ram_width = 19;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 4;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 15;
defparam ram_block1a16.port_b_logical_ram_depth = 16;
defparam ram_block1a16.port_b_logical_ram_width = 19;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 4;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 15;
defparam ram_block1a17.port_a_logical_ram_depth = 16;
defparam ram_block1a17.port_a_logical_ram_width = 19;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 4;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 15;
defparam ram_block1a17.port_b_logical_ram_depth = 16;
defparam ram_block1a17.port_b_logical_ram_width = 19;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[2].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 4;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 15;
defparam ram_block1a18.port_a_logical_ram_depth = 16;
defparam ram_block1a18.port_a_logical_ram_width = 19;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 4;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 15;
defparam ram_block1a18.port_b_logical_ram_depth = 16;
defparam ram_block1a18.port_b_logical_ram_width = 19;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

endmodule

module cic_cntr_ika_2 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout());
defparam counter_comb_bita2.lut_mask = 16'h5A5A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

endmodule

module cic_cntr_jka_2 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module cic_cntr_vk6_2 (
	full_dff,
	counter_reg_bit_1,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_0,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_1;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_0;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_channel_buffer_3 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_3,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_3;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_4 buffer_FIFO(
	.q({q_unconnected_wire_22,q_unconnected_wire_21,q_unconnected_wire_20,q_unconnected_wire_19,q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({gnd,gnd,gnd,gnd,data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_3(fifo_rdreq_3),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module cic_scfifo_4 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_3,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[22:0] q;
input 	[22:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_3;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_1351_3 auto_generated(
	.q({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_3(fifo_rdreq_3),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module cic_scfifo_1351_3 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_3,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_3;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_a_dpfifo_c0u_3 dpfifo(
	.q({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_3(fifo_rdreq_3),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module cic_a_dpfifo_c0u_3 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_3,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_3;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \empty_dff~2_combout ;


cic_cntr_jka_3 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_cntr_vk6_3 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_cntr_ika_3 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_altsyncram_dlg1_3 FIFOram(
	.q_b({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data_a({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock0(clock),
	.clock1(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

fiftyfivenm_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

fiftyfivenm_lcell_comb \valid_rreq~0 (
	.dataa(fifo_rdreq_3),
	.datab(\empty_dff~q ),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(\usedw_counter|counter_reg_bit[3]~q ),
	.datac(\usedw_counter|counter_reg_bit[2]~q ),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hFEFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \_~1 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~0_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFEFF;
defparam \_~1 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

fiftyfivenm_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(\usedw_counter|counter_reg_bit[0]~q ),
	.datac(\usedw_counter|counter_reg_bit[3]~q ),
	.datad(\usedw_counter|counter_reg_bit[2]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~2 (
	.dataa(stall_reg),
	.datab(fifo_rdreq_3),
	.datac(\empty_dff~q ),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFFFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~1 (
	.dataa(fifo_rdreq_3),
	.datab(\empty_dff~q ),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

endmodule

module cic_altsyncram_dlg1_3 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q_b;
input 	[18:0] data_a;
input 	[3:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[3:0] address_b;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

fiftyfivenm_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk1_output_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 19;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 19;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk1_output_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 19;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 19;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk1_output_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 19;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 19;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk1_output_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 19;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 19;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk1_output_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 19;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 19;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 19;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 19;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 19;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 19;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 19;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 19;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 19;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 19;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 19;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 19;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 19;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 19;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 19;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 19;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 19;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 19;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 19;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 19;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 19;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 19;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 19;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 19;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 4;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 15;
defparam ram_block1a16.port_a_logical_ram_depth = 16;
defparam ram_block1a16.port_a_logical_ram_width = 19;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 4;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 15;
defparam ram_block1a16.port_b_logical_ram_depth = 16;
defparam ram_block1a16.port_b_logical_ram_width = 19;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 4;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 15;
defparam ram_block1a17.port_a_logical_ram_depth = 16;
defparam ram_block1a17.port_a_logical_ram_width = 19;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 4;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 15;
defparam ram_block1a17.port_b_logical_ram_depth = 16;
defparam ram_block1a17.port_b_logical_ram_width = 19;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[3].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 4;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 15;
defparam ram_block1a18.port_a_logical_ram_depth = 16;
defparam ram_block1a18.port_a_logical_ram_width = 19;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 4;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 15;
defparam ram_block1a18.port_b_logical_ram_depth = 16;
defparam ram_block1a18.port_b_logical_ram_width = 19;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

endmodule

module cic_cntr_ika_3 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout());
defparam counter_comb_bita2.lut_mask = 16'h5A5A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

endmodule

module cic_cntr_jka_3 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module cic_cntr_vk6_3 (
	full_dff,
	counter_reg_bit_1,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_0,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_1;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_0;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_channel_buffer_4 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_4,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_4;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_5 buffer_FIFO(
	.q({q_unconnected_wire_22,q_unconnected_wire_21,q_unconnected_wire_20,q_unconnected_wire_19,q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({gnd,gnd,gnd,gnd,data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_4(fifo_rdreq_4),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module cic_scfifo_5 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_4,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[22:0] q;
input 	[22:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_4;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_1351_4 auto_generated(
	.q({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_4(fifo_rdreq_4),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module cic_scfifo_1351_4 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_4,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_4;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_a_dpfifo_c0u_4 dpfifo(
	.q({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_4(fifo_rdreq_4),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module cic_a_dpfifo_c0u_4 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_4,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_4;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \empty_dff~2_combout ;


cic_cntr_jka_4 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_cntr_vk6_4 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_cntr_ika_4 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_altsyncram_dlg1_4 FIFOram(
	.q_b({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data_a({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock0(clock),
	.clock1(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

fiftyfivenm_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

fiftyfivenm_lcell_comb \valid_rreq~0 (
	.dataa(fifo_rdreq_4),
	.datab(\empty_dff~q ),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(\usedw_counter|counter_reg_bit[3]~q ),
	.datac(\usedw_counter|counter_reg_bit[2]~q ),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hFEFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \_~1 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~0_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFEFF;
defparam \_~1 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

fiftyfivenm_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(\usedw_counter|counter_reg_bit[0]~q ),
	.datac(\usedw_counter|counter_reg_bit[3]~q ),
	.datad(\usedw_counter|counter_reg_bit[2]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~2 (
	.dataa(stall_reg),
	.datab(fifo_rdreq_4),
	.datac(\empty_dff~q ),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFFFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~1 (
	.dataa(fifo_rdreq_4),
	.datab(\empty_dff~q ),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

endmodule

module cic_altsyncram_dlg1_4 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q_b;
input 	[18:0] data_a;
input 	[3:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[3:0] address_b;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

fiftyfivenm_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk1_output_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 19;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 19;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk1_output_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 19;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 19;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk1_output_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 19;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 19;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk1_output_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 19;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 19;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk1_output_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 19;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 19;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 19;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 19;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 19;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 19;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 19;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 19;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 19;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 19;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 19;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 19;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 19;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 19;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 19;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 19;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 19;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 19;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 19;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 19;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 19;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 19;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 19;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 19;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 4;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 15;
defparam ram_block1a16.port_a_logical_ram_depth = 16;
defparam ram_block1a16.port_a_logical_ram_width = 19;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 4;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 15;
defparam ram_block1a16.port_b_logical_ram_depth = 16;
defparam ram_block1a16.port_b_logical_ram_width = 19;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 4;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 15;
defparam ram_block1a17.port_a_logical_ram_depth = 16;
defparam ram_block1a17.port_a_logical_ram_width = 19;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 4;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 15;
defparam ram_block1a17.port_b_logical_ram_depth = 16;
defparam ram_block1a17.port_b_logical_ram_width = 19;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[4].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 4;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 15;
defparam ram_block1a18.port_a_logical_ram_depth = 16;
defparam ram_block1a18.port_a_logical_ram_width = 19;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 4;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 15;
defparam ram_block1a18.port_b_logical_ram_depth = 16;
defparam ram_block1a18.port_b_logical_ram_width = 19;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

endmodule

module cic_cntr_ika_4 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout());
defparam counter_comb_bita2.lut_mask = 16'h5A5A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

endmodule

module cic_cntr_jka_4 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module cic_cntr_vk6_4 (
	full_dff,
	counter_reg_bit_1,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_0,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_1;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_0;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_channel_buffer_5 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_5,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_5;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_6 buffer_FIFO(
	.q({q_unconnected_wire_22,q_unconnected_wire_21,q_unconnected_wire_20,q_unconnected_wire_19,q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({gnd,gnd,gnd,gnd,data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_5(fifo_rdreq_5),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module cic_scfifo_6 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_5,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[22:0] q;
input 	[22:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_5;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_1351_5 auto_generated(
	.q({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_5(fifo_rdreq_5),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module cic_scfifo_1351_5 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_5,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_5;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_a_dpfifo_c0u_5 dpfifo(
	.q({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_5(fifo_rdreq_5),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module cic_a_dpfifo_c0u_5 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_5,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_5;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \empty_dff~2_combout ;


cic_cntr_jka_5 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_cntr_vk6_5 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_cntr_ika_5 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_altsyncram_dlg1_5 FIFOram(
	.q_b({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data_a({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock0(clock),
	.clock1(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

fiftyfivenm_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

fiftyfivenm_lcell_comb \valid_rreq~0 (
	.dataa(fifo_rdreq_5),
	.datab(\empty_dff~q ),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(\usedw_counter|counter_reg_bit[3]~q ),
	.datac(\usedw_counter|counter_reg_bit[2]~q ),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hFEFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \_~1 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~0_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFEFF;
defparam \_~1 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

fiftyfivenm_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~0 (
	.dataa(valid_wreq),
	.datab(\full_dff~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(\usedw_counter|counter_reg_bit[0]~q ),
	.datac(\usedw_counter|counter_reg_bit[3]~q ),
	.datad(\usedw_counter|counter_reg_bit[2]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~2 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~1_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~0_combout ),
	.datac(\usedw_will_be_1~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFEFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~1 (
	.dataa(fifo_rdreq_5),
	.datab(\empty_dff~q ),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

endmodule

module cic_altsyncram_dlg1_5 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q_b;
input 	[18:0] data_a;
input 	[3:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[3:0] address_b;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

fiftyfivenm_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk1_output_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 19;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 19;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk1_output_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 19;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 19;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk1_output_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 19;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 19;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk1_output_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 19;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 19;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk1_output_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 19;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 19;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 19;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 19;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 19;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 19;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 19;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 19;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 19;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 19;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 19;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 19;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 19;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 19;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 19;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 19;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 19;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 19;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 19;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 19;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 19;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 19;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 19;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 19;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 4;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 15;
defparam ram_block1a16.port_a_logical_ram_depth = 16;
defparam ram_block1a16.port_a_logical_ram_width = 19;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 4;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 15;
defparam ram_block1a16.port_b_logical_ram_depth = 16;
defparam ram_block1a16.port_b_logical_ram_width = 19;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 4;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 15;
defparam ram_block1a17.port_a_logical_ram_depth = 16;
defparam ram_block1a17.port_a_logical_ram_width = 19;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 4;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 15;
defparam ram_block1a17.port_b_logical_ram_depth = 16;
defparam ram_block1a17.port_b_logical_ram_width = 19;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[5].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 4;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 15;
defparam ram_block1a18.port_a_logical_ram_depth = 16;
defparam ram_block1a18.port_a_logical_ram_width = 19;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 4;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 15;
defparam ram_block1a18.port_b_logical_ram_depth = 16;
defparam ram_block1a18.port_b_logical_ram_width = 19;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

endmodule

module cic_cntr_ika_5 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout());
defparam counter_comb_bita2.lut_mask = 16'h5A5A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

endmodule

module cic_cntr_jka_5 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module cic_cntr_vk6_5 (
	full_dff,
	counter_reg_bit_1,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_0,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_1;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_0;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_channel_buffer_6 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_6,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_6;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_7 buffer_FIFO(
	.q({q_unconnected_wire_22,q_unconnected_wire_21,q_unconnected_wire_20,q_unconnected_wire_19,q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({gnd,gnd,gnd,gnd,data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_6(fifo_rdreq_6),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module cic_scfifo_7 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_6,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[22:0] q;
input 	[22:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_6;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_1351_6 auto_generated(
	.q({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_6(fifo_rdreq_6),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module cic_scfifo_1351_6 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_6,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_6;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_a_dpfifo_c0u_6 dpfifo(
	.q({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_6(fifo_rdreq_6),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module cic_a_dpfifo_c0u_6 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_6,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_6;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \empty_dff~2_combout ;
wire \usedw_will_be_1~3_combout ;


cic_cntr_jka_6 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_cntr_vk6_6 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_cntr_ika_6 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_altsyncram_dlg1_6 FIFOram(
	.q_b({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data_a({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock0(clock),
	.clock1(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

fiftyfivenm_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

fiftyfivenm_lcell_comb \valid_rreq~0 (
	.dataa(fifo_rdreq_6),
	.datab(\empty_dff~q ),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(\usedw_counter|counter_reg_bit[3]~q ),
	.datac(\usedw_counter|counter_reg_bit[2]~q ),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hFEFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \_~1 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~0_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFEFF;
defparam \_~1 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

fiftyfivenm_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(\usedw_counter|counter_reg_bit[0]~q ),
	.datac(\usedw_counter|counter_reg_bit[3]~q ),
	.datad(\usedw_counter|counter_reg_bit[2]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~2 (
	.dataa(\usedw_will_be_1~1_combout ),
	.datab(\valid_wreq~0_combout ),
	.datac(\valid_rreq~0_combout ),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hEFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~1 (
	.dataa(fifo_rdreq_6),
	.datab(\empty_dff~q ),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hEEEE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

endmodule

module cic_altsyncram_dlg1_6 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q_b;
input 	[18:0] data_a;
input 	[3:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[3:0] address_b;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

fiftyfivenm_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk1_output_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 19;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 19;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk1_output_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 19;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 19;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk1_output_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 19;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 19;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk1_output_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 19;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 19;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk1_output_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 19;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 19;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 19;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 19;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 19;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 19;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 19;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 19;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 19;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 19;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 19;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 19;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 19;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 19;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 19;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 19;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 19;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 19;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 19;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 19;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 19;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 19;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 19;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 19;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 4;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 15;
defparam ram_block1a16.port_a_logical_ram_depth = 16;
defparam ram_block1a16.port_a_logical_ram_width = 19;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 4;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 15;
defparam ram_block1a16.port_b_logical_ram_depth = 16;
defparam ram_block1a16.port_b_logical_ram_width = 19;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 4;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 15;
defparam ram_block1a17.port_a_logical_ram_depth = 16;
defparam ram_block1a17.port_a_logical_ram_width = 19;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 4;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 15;
defparam ram_block1a17.port_b_logical_ram_depth = 16;
defparam ram_block1a17.port_b_logical_ram_width = 19;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[6].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 4;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 15;
defparam ram_block1a18.port_a_logical_ram_depth = 16;
defparam ram_block1a18.port_a_logical_ram_width = 19;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 4;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 15;
defparam ram_block1a18.port_b_logical_ram_depth = 16;
defparam ram_block1a18.port_b_logical_ram_width = 19;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

endmodule

module cic_cntr_ika_6 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout());
defparam counter_comb_bita2.lut_mask = 16'h5A5A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

endmodule

module cic_cntr_jka_6 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module cic_cntr_vk6_6 (
	full_dff,
	counter_reg_bit_1,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_0,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_1;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_0;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_channel_buffer_7 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_7,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_7;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_8 buffer_FIFO(
	.q({q_unconnected_wire_22,q_unconnected_wire_21,q_unconnected_wire_20,q_unconnected_wire_19,q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({gnd,gnd,gnd,gnd,data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_7(fifo_rdreq_7),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module cic_scfifo_8 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_7,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[22:0] q;
input 	[22:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_7;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_1351_7 auto_generated(
	.q({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_7(fifo_rdreq_7),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module cic_scfifo_1351_7 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_7,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_7;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_a_dpfifo_c0u_7 dpfifo(
	.q({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_7(fifo_rdreq_7),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module cic_a_dpfifo_c0u_7 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_7,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_7;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \empty_dff~2_combout ;


cic_cntr_jka_7 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_cntr_vk6_7 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_cntr_ika_7 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_altsyncram_dlg1_7 FIFOram(
	.q_b({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data_a({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock0(clock),
	.clock1(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

fiftyfivenm_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

fiftyfivenm_lcell_comb \valid_rreq~0 (
	.dataa(fifo_rdreq_7),
	.datab(\empty_dff~q ),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(\usedw_counter|counter_reg_bit[3]~q ),
	.datac(\usedw_counter|counter_reg_bit[2]~q ),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hFEFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \_~1 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~0_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFEFF;
defparam \_~1 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

fiftyfivenm_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~0 (
	.dataa(valid_wreq),
	.datab(\full_dff~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(\usedw_counter|counter_reg_bit[0]~q ),
	.datac(\usedw_counter|counter_reg_bit[3]~q ),
	.datad(\usedw_counter|counter_reg_bit[2]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~2 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~1_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~0_combout ),
	.datac(\usedw_will_be_1~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFEFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~1 (
	.dataa(fifo_rdreq_7),
	.datab(\empty_dff~q ),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

endmodule

module cic_altsyncram_dlg1_7 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q_b;
input 	[18:0] data_a;
input 	[3:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[3:0] address_b;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

fiftyfivenm_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk1_output_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 19;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 19;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk1_output_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 19;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 19;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk1_output_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 19;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 19;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk1_output_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 19;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 19;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk1_output_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 19;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 19;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 19;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 19;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 19;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 19;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 19;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 19;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 19;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 19;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 19;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 19;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 19;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 19;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 19;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 19;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 19;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 19;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 19;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 19;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 19;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 19;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 19;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 19;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 4;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 15;
defparam ram_block1a16.port_a_logical_ram_depth = 16;
defparam ram_block1a16.port_a_logical_ram_width = 19;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 4;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 15;
defparam ram_block1a16.port_b_logical_ram_depth = 16;
defparam ram_block1a16.port_b_logical_ram_width = 19;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 4;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 15;
defparam ram_block1a17.port_a_logical_ram_depth = 16;
defparam ram_block1a17.port_a_logical_ram_width = 19;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 4;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 15;
defparam ram_block1a17.port_b_logical_ram_depth = 16;
defparam ram_block1a17.port_b_logical_ram_width = 19;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[7].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 4;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 15;
defparam ram_block1a18.port_a_logical_ram_depth = 16;
defparam ram_block1a18.port_a_logical_ram_width = 19;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 4;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 15;
defparam ram_block1a18.port_b_logical_ram_depth = 16;
defparam ram_block1a18.port_b_logical_ram_width = 19;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

endmodule

module cic_cntr_ika_7 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout());
defparam counter_comb_bita2.lut_mask = 16'h5A5A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

endmodule

module cic_cntr_jka_7 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module cic_cntr_vk6_7 (
	full_dff,
	counter_reg_bit_1,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_0,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_1;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_0;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_channel_buffer_8 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_8,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_8;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_9 buffer_FIFO(
	.q({q_unconnected_wire_22,q_unconnected_wire_21,q_unconnected_wire_20,q_unconnected_wire_19,q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({gnd,gnd,gnd,gnd,data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_8(fifo_rdreq_8),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module cic_scfifo_9 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_8,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[22:0] q;
input 	[22:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_8;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_1351_8 auto_generated(
	.q({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_8(fifo_rdreq_8),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module cic_scfifo_1351_8 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_8,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_8;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_a_dpfifo_c0u_8 dpfifo(
	.q({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.valid_wreq(valid_wreq),
	.fifo_rdreq_8(fifo_rdreq_8),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module cic_a_dpfifo_c0u_8 (
	q,
	data,
	stall_reg,
	valid_wreq,
	fifo_rdreq_8,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q;
input 	[18:0] data;
input 	stall_reg;
input 	valid_wreq;
input 	fifo_rdreq_8;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \full_dff~q ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[1]~q ;
wire \usedw_counter|counter_reg_bit[3]~q ;
wire \usedw_counter|counter_reg_bit[2]~q ;
wire \usedw_counter|counter_reg_bit[0]~q ;
wire \valid_wreq~0_combout ;
wire \empty_dff~q ;
wire \valid_rreq~0_combout ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \_~0_combout ;
wire \_~1_combout ;
wire \usedw_is_0_dff~q ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \empty_dff~1_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \empty_dff~2_combout ;


cic_cntr_jka_8 wr_ptr(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.valid_wreq(valid_wreq),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_cntr_vk6_8 usedw_counter(
	.full_dff(\full_dff~q ),
	.counter_reg_bit_1(\usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_3(\usedw_counter|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_0(\usedw_counter|counter_reg_bit[0]~q ),
	.valid_wreq(valid_wreq),
	.updown(\valid_wreq~0_combout ),
	.valid_rreq(\valid_rreq~0_combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_cntr_ika_8 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.valid_rreq(\valid_rreq~0_combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_altsyncram_dlg1_8 FIFOram(
	.q_b({q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data_a({data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~0_combout ),
	.clocken1(\valid_rreq~0_combout ),
	.address_b({\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock0(clock),
	.clock1(clock));

dffeas full_dff(
	.clk(clock),
	.d(\_~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

fiftyfivenm_lcell_comb \valid_wreq~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(gnd),
	.datad(\full_dff~q ),
	.cin(gnd),
	.combout(\valid_wreq~0_combout ),
	.cout());
defparam \valid_wreq~0 .lut_mask = 16'hAAFF;
defparam \valid_wreq~0 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

fiftyfivenm_lcell_comb \valid_rreq~0 (
	.dataa(fifo_rdreq_8),
	.datab(\empty_dff~q ),
	.datac(gnd),
	.datad(stall_reg),
	.cin(gnd),
	.combout(\valid_rreq~0_combout ),
	.cout());
defparam \valid_rreq~0 .lut_mask = 16'hEEFF;
defparam \valid_rreq~0 .sum_lutc_input = "datac";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(\usedw_counter|counter_reg_bit[3]~q ),
	.datac(\usedw_counter|counter_reg_bit[2]~q ),
	.datad(\usedw_counter|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hFEFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \_~1 (
	.dataa(\full_dff~q ),
	.datab(valid_wreq),
	.datac(\_~0_combout ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hFEFF;
defparam \_~1 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

fiftyfivenm_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~0_combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~0 (
	.dataa(\usedw_counter|counter_reg_bit[1]~q ),
	.datab(\usedw_counter|counter_reg_bit[0]~q ),
	.datac(\usedw_counter|counter_reg_bit[3]~q ),
	.datad(\usedw_counter|counter_reg_bit[2]~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~0_combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~2 (
	.dataa(stall_reg),
	.datab(fifo_rdreq_8),
	.datac(\empty_dff~q ),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~2_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFFFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~0_combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~0_combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~1 (
	.dataa(fifo_rdreq_8),
	.datab(\empty_dff~q ),
	.datac(stall_reg),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(\valid_rreq~0_combout ),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

endmodule

module cic_altsyncram_dlg1_8 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[18:0] q_b;
input 	[18:0] data_a;
input 	[3:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[3:0] address_b;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

fiftyfivenm_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk1_output_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 19;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 4;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 15;
defparam ram_block1a0.port_b_logical_ram_depth = 16;
defparam ram_block1a0.port_b_logical_ram_width = 19;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk1_output_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 19;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 4;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 15;
defparam ram_block1a1.port_b_logical_ram_depth = 16;
defparam ram_block1a1.port_b_logical_ram_width = 19;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk1_output_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 19;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 4;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 15;
defparam ram_block1a2.port_b_logical_ram_depth = 16;
defparam ram_block1a2.port_b_logical_ram_width = 19;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk1_output_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 19;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 4;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 15;
defparam ram_block1a3.port_b_logical_ram_depth = 16;
defparam ram_block1a3.port_b_logical_ram_width = 19;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk1_output_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 19;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 4;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 15;
defparam ram_block1a4.port_b_logical_ram_depth = 16;
defparam ram_block1a4.port_b_logical_ram_width = 19;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 19;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 4;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 15;
defparam ram_block1a5.port_b_logical_ram_depth = 16;
defparam ram_block1a5.port_b_logical_ram_width = 19;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 19;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 4;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 15;
defparam ram_block1a6.port_b_logical_ram_depth = 16;
defparam ram_block1a6.port_b_logical_ram_width = 19;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 19;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 4;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 15;
defparam ram_block1a7.port_b_logical_ram_depth = 16;
defparam ram_block1a7.port_b_logical_ram_width = 19;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 19;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 4;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 15;
defparam ram_block1a8.port_b_logical_ram_depth = 16;
defparam ram_block1a8.port_b_logical_ram_width = 19;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 19;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 4;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 15;
defparam ram_block1a9.port_b_logical_ram_depth = 16;
defparam ram_block1a9.port_b_logical_ram_width = 19;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 19;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 4;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 15;
defparam ram_block1a10.port_b_logical_ram_depth = 16;
defparam ram_block1a10.port_b_logical_ram_width = 19;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 19;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 4;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 15;
defparam ram_block1a11.port_b_logical_ram_depth = 16;
defparam ram_block1a11.port_b_logical_ram_width = 19;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 19;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 4;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 15;
defparam ram_block1a12.port_b_logical_ram_depth = 16;
defparam ram_block1a12.port_b_logical_ram_width = 19;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 19;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 4;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 15;
defparam ram_block1a13.port_b_logical_ram_depth = 16;
defparam ram_block1a13.port_b_logical_ram_width = 19;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 19;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 4;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 15;
defparam ram_block1a14.port_b_logical_ram_depth = 16;
defparam ram_block1a14.port_b_logical_ram_width = 19;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 19;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 4;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 15;
defparam ram_block1a15.port_b_logical_ram_depth = 16;
defparam ram_block1a15.port_b_logical_ram_width = 19;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 4;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 15;
defparam ram_block1a16.port_a_logical_ram_depth = 16;
defparam ram_block1a16.port_a_logical_ram_width = 19;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 4;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 15;
defparam ram_block1a16.port_b_logical_ram_depth = 16;
defparam ram_block1a16.port_b_logical_ram_width = 19;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 4;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 15;
defparam ram_block1a17.port_a_logical_ram_depth = 16;
defparam ram_block1a17.port_a_logical_ram_width = 19;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 4;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 15;
defparam ram_block1a17.port_b_logical_ram_depth = 16;
defparam ram_block1a17.port_b_logical_ram_width = 19;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_channel_buffer:integrator[8].fifo_regulator|scfifo:buffer_FIFO|scfifo_1351:auto_generated|a_dpfifo_c0u:dpfifo|altsyncram_dlg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 4;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 15;
defparam ram_block1a18.port_a_logical_ram_depth = 16;
defparam ram_block1a18.port_a_logical_ram_width = 19;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 4;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 15;
defparam ram_block1a18.port_b_logical_ram_depth = 16;
defparam ram_block1a18.port_b_logical_ram_width = 19;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

endmodule

module cic_cntr_ika_8 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout());
defparam counter_comb_bita2.lut_mask = 16'h5A5A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

endmodule

module cic_cntr_jka_8 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_wreq),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module cic_cntr_vk6_8 (
	full_dff,
	counter_reg_bit_1,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_0,
	valid_wreq,
	updown,
	valid_rreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_1;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_0;
input 	valid_wreq;
input 	updown;
input 	valid_rreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \_~0_combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(full_dff),
	.datac(valid_wreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h96FF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_differentiator (
	dout_0,
	dout_1,
	dout_2,
	dout_3,
	dout_4,
	dout_5,
	dout_6,
	dout_7,
	dout_8,
	dout_9,
	dout_10,
	dout_11,
	dout_12,
	dout_13,
	dout_14,
	dout_15,
	dout_16,
	dout_17,
	dout_18,
	stall_reg,
	ena_diff_s_1,
	dout_valid1,
	ena_diff_s_11,
	Mux18,
	Mux14,
	Mux13,
	Mux12,
	Mux11,
	Mux10,
	Mux9,
	Mux8,
	Mux7,
	Mux6,
	Mux5,
	Mux4,
	Mux3,
	Mux2,
	Mux1,
	Mux0,
	Mux17,
	Mux16,
	Mux15,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dout_0;
output 	dout_1;
output 	dout_2;
output 	dout_3;
output 	dout_4;
output 	dout_5;
output 	dout_6;
output 	dout_7;
output 	dout_8;
output 	dout_9;
output 	dout_10;
output 	dout_11;
output 	dout_12;
output 	dout_13;
output 	dout_14;
output 	dout_15;
output 	dout_16;
output 	dout_17;
output 	dout_18;
input 	stall_reg;
input 	ena_diff_s_1;
output 	dout_valid1;
input 	ena_diff_s_11;
input 	Mux18;
input 	Mux14;
input 	Mux13;
input 	Mux12;
input 	Mux11;
input 	Mux10;
input 	Mux9;
input 	Mux8;
input 	Mux7;
input 	Mux6;
input 	Mux5;
input 	Mux4;
input 	Mux3;
input 	Mux2;
input 	Mux1;
input 	Mux0;
input 	Mux17;
input 	Mux16;
input 	Mux15;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0~portbdataout ;
wire \ena_and_valid~combout ;
wire \dout[0]~19_combout ;
wire \dout[8]~21_combout ;
wire \dout[0]~20 ;
wire \dout[1]~22_combout ;
wire \dout[1]~23 ;
wire \dout[2]~24_combout ;
wire \dout[2]~25 ;
wire \dout[3]~26_combout ;
wire \dout[3]~27 ;
wire \dout[4]~28_combout ;
wire \dout[4]~29 ;
wire \dout[5]~30_combout ;
wire \dout[5]~31 ;
wire \dout[6]~32_combout ;
wire \dout[6]~33 ;
wire \dout[7]~34_combout ;
wire \dout[7]~35 ;
wire \dout[8]~36_combout ;
wire \dout[8]~37 ;
wire \dout[9]~38_combout ;
wire \dout[9]~39 ;
wire \dout[10]~40_combout ;
wire \dout[10]~41 ;
wire \dout[11]~42_combout ;
wire \dout[11]~43 ;
wire \dout[12]~44_combout ;
wire \dout[12]~45 ;
wire \dout[13]~46_combout ;
wire \dout[13]~47 ;
wire \dout[14]~48_combout ;
wire \dout[14]~49 ;
wire \dout[15]~50_combout ;
wire \dout[15]~51 ;
wire \dout[16]~52_combout ;
wire \dout[16]~53 ;
wire \dout[17]~54_combout ;
wire \dout[17]~55 ;
wire \dout[18]~56_combout ;
wire \dout_valid~0_combout ;


cic_auk_dspip_delay \glogic:u0 (
	.ram_block5a18(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18~portbdataout ),
	.ram_block5a17(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17~portbdataout ),
	.ram_block5a16(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16~portbdataout ),
	.ram_block5a15(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15~portbdataout ),
	.ram_block5a14(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14~portbdataout ),
	.ram_block5a13(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13~portbdataout ),
	.ram_block5a12(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12~portbdataout ),
	.ram_block5a11(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11~portbdataout ),
	.ram_block5a10(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10~portbdataout ),
	.ram_block5a9(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9~portbdataout ),
	.ram_block5a8(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8~portbdataout ),
	.ram_block5a7(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7~portbdataout ),
	.ram_block5a6(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6~portbdataout ),
	.ram_block5a5(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5~portbdataout ),
	.ram_block5a4(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4~portbdataout ),
	.ram_block5a3(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3~portbdataout ),
	.ram_block5a2(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2~portbdataout ),
	.ram_block5a1(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1~portbdataout ),
	.ram_block5a0(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0~portbdataout ),
	.stall_reg(stall_reg),
	.ena_diff_s_1(ena_diff_s_11),
	.Mux18(Mux18),
	.Mux14(Mux14),
	.Mux13(Mux13),
	.Mux12(Mux12),
	.Mux11(Mux11),
	.Mux10(Mux10),
	.Mux9(Mux9),
	.Mux8(Mux8),
	.Mux7(Mux7),
	.Mux6(Mux6),
	.Mux5(Mux5),
	.Mux4(Mux4),
	.Mux3(Mux3),
	.Mux2(Mux2),
	.Mux1(Mux1),
	.Mux0(Mux0),
	.ena_and_valid(\ena_and_valid~combout ),
	.Mux17(Mux17),
	.Mux16(Mux16),
	.Mux15(Mux15),
	.clk(clk),
	.reset_n(reset_n));

fiftyfivenm_lcell_comb ena_and_valid(
	.dataa(stall_reg),
	.datab(gnd),
	.datac(gnd),
	.datad(ena_diff_s_11),
	.cin(gnd),
	.combout(\ena_and_valid~combout ),
	.cout());
defparam ena_and_valid.lut_mask = 16'hFF55;
defparam ena_and_valid.sum_lutc_input = "datac";

dffeas \dout[0] (
	.clk(clk),
	.d(\dout[0]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[8]~21_combout ),
	.q(dout_0),
	.prn(vcc));
defparam \dout[0] .is_wysiwyg = "true";
defparam \dout[0] .power_up = "low";

dffeas \dout[1] (
	.clk(clk),
	.d(\dout[1]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[8]~21_combout ),
	.q(dout_1),
	.prn(vcc));
defparam \dout[1] .is_wysiwyg = "true";
defparam \dout[1] .power_up = "low";

dffeas \dout[2] (
	.clk(clk),
	.d(\dout[2]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[8]~21_combout ),
	.q(dout_2),
	.prn(vcc));
defparam \dout[2] .is_wysiwyg = "true";
defparam \dout[2] .power_up = "low";

dffeas \dout[3] (
	.clk(clk),
	.d(\dout[3]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[8]~21_combout ),
	.q(dout_3),
	.prn(vcc));
defparam \dout[3] .is_wysiwyg = "true";
defparam \dout[3] .power_up = "low";

dffeas \dout[4] (
	.clk(clk),
	.d(\dout[4]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[8]~21_combout ),
	.q(dout_4),
	.prn(vcc));
defparam \dout[4] .is_wysiwyg = "true";
defparam \dout[4] .power_up = "low";

dffeas \dout[5] (
	.clk(clk),
	.d(\dout[5]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[8]~21_combout ),
	.q(dout_5),
	.prn(vcc));
defparam \dout[5] .is_wysiwyg = "true";
defparam \dout[5] .power_up = "low";

dffeas \dout[6] (
	.clk(clk),
	.d(\dout[6]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[8]~21_combout ),
	.q(dout_6),
	.prn(vcc));
defparam \dout[6] .is_wysiwyg = "true";
defparam \dout[6] .power_up = "low";

dffeas \dout[7] (
	.clk(clk),
	.d(\dout[7]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[8]~21_combout ),
	.q(dout_7),
	.prn(vcc));
defparam \dout[7] .is_wysiwyg = "true";
defparam \dout[7] .power_up = "low";

dffeas \dout[8] (
	.clk(clk),
	.d(\dout[8]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[8]~21_combout ),
	.q(dout_8),
	.prn(vcc));
defparam \dout[8] .is_wysiwyg = "true";
defparam \dout[8] .power_up = "low";

dffeas \dout[9] (
	.clk(clk),
	.d(\dout[9]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[8]~21_combout ),
	.q(dout_9),
	.prn(vcc));
defparam \dout[9] .is_wysiwyg = "true";
defparam \dout[9] .power_up = "low";

dffeas \dout[10] (
	.clk(clk),
	.d(\dout[10]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[8]~21_combout ),
	.q(dout_10),
	.prn(vcc));
defparam \dout[10] .is_wysiwyg = "true";
defparam \dout[10] .power_up = "low";

dffeas \dout[11] (
	.clk(clk),
	.d(\dout[11]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[8]~21_combout ),
	.q(dout_11),
	.prn(vcc));
defparam \dout[11] .is_wysiwyg = "true";
defparam \dout[11] .power_up = "low";

dffeas \dout[12] (
	.clk(clk),
	.d(\dout[12]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[8]~21_combout ),
	.q(dout_12),
	.prn(vcc));
defparam \dout[12] .is_wysiwyg = "true";
defparam \dout[12] .power_up = "low";

dffeas \dout[13] (
	.clk(clk),
	.d(\dout[13]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[8]~21_combout ),
	.q(dout_13),
	.prn(vcc));
defparam \dout[13] .is_wysiwyg = "true";
defparam \dout[13] .power_up = "low";

dffeas \dout[14] (
	.clk(clk),
	.d(\dout[14]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[8]~21_combout ),
	.q(dout_14),
	.prn(vcc));
defparam \dout[14] .is_wysiwyg = "true";
defparam \dout[14] .power_up = "low";

dffeas \dout[15] (
	.clk(clk),
	.d(\dout[15]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[8]~21_combout ),
	.q(dout_15),
	.prn(vcc));
defparam \dout[15] .is_wysiwyg = "true";
defparam \dout[15] .power_up = "low";

dffeas \dout[16] (
	.clk(clk),
	.d(\dout[16]~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[8]~21_combout ),
	.q(dout_16),
	.prn(vcc));
defparam \dout[16] .is_wysiwyg = "true";
defparam \dout[16] .power_up = "low";

dffeas \dout[17] (
	.clk(clk),
	.d(\dout[17]~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[8]~21_combout ),
	.q(dout_17),
	.prn(vcc));
defparam \dout[17] .is_wysiwyg = "true";
defparam \dout[17] .power_up = "low";

dffeas \dout[18] (
	.clk(clk),
	.d(\dout[18]~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[8]~21_combout ),
	.q(dout_18),
	.prn(vcc));
defparam \dout[18] .is_wysiwyg = "true";
defparam \dout[18] .power_up = "low";

dffeas dout_valid(
	.clk(clk),
	.d(\dout_valid~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena_diff_s_1),
	.q(dout_valid1),
	.prn(vcc));
defparam dout_valid.is_wysiwyg = "true";
defparam dout_valid.power_up = "low";

fiftyfivenm_lcell_comb \dout[0]~19 (
	.dataa(Mux18),
	.datab(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18~portbdataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\dout[0]~19_combout ),
	.cout(\dout[0]~20 ));
defparam \dout[0]~19 .lut_mask = 16'h66BB;
defparam \dout[0]~19 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dout[8]~21 (
	.dataa(reset_n),
	.datab(stall_reg),
	.datac(gnd),
	.datad(ena_diff_s_11),
	.cin(gnd),
	.combout(\dout[8]~21_combout ),
	.cout());
defparam \dout[8]~21 .lut_mask = 16'hFF77;
defparam \dout[8]~21 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dout[1]~22 (
	.dataa(Mux17),
	.datab(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17~portbdataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[0]~20 ),
	.combout(\dout[1]~22_combout ),
	.cout(\dout[1]~23 ));
defparam \dout[1]~22 .lut_mask = 16'h96DF;
defparam \dout[1]~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[2]~24 (
	.dataa(Mux16),
	.datab(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16~portbdataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[1]~23 ),
	.combout(\dout[2]~24_combout ),
	.cout(\dout[2]~25 ));
defparam \dout[2]~24 .lut_mask = 16'h96BF;
defparam \dout[2]~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[3]~26 (
	.dataa(Mux15),
	.datab(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15~portbdataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[2]~25 ),
	.combout(\dout[3]~26_combout ),
	.cout(\dout[3]~27 ));
defparam \dout[3]~26 .lut_mask = 16'h96DF;
defparam \dout[3]~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[4]~28 (
	.dataa(Mux14),
	.datab(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14~portbdataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[3]~27 ),
	.combout(\dout[4]~28_combout ),
	.cout(\dout[4]~29 ));
defparam \dout[4]~28 .lut_mask = 16'h96BF;
defparam \dout[4]~28 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[5]~30 (
	.dataa(Mux13),
	.datab(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13~portbdataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[4]~29 ),
	.combout(\dout[5]~30_combout ),
	.cout(\dout[5]~31 ));
defparam \dout[5]~30 .lut_mask = 16'h96DF;
defparam \dout[5]~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[6]~32 (
	.dataa(Mux12),
	.datab(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12~portbdataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[5]~31 ),
	.combout(\dout[6]~32_combout ),
	.cout(\dout[6]~33 ));
defparam \dout[6]~32 .lut_mask = 16'h96BF;
defparam \dout[6]~32 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[7]~34 (
	.dataa(Mux11),
	.datab(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11~portbdataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[6]~33 ),
	.combout(\dout[7]~34_combout ),
	.cout(\dout[7]~35 ));
defparam \dout[7]~34 .lut_mask = 16'h96DF;
defparam \dout[7]~34 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[8]~36 (
	.dataa(Mux10),
	.datab(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10~portbdataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[7]~35 ),
	.combout(\dout[8]~36_combout ),
	.cout(\dout[8]~37 ));
defparam \dout[8]~36 .lut_mask = 16'h96BF;
defparam \dout[8]~36 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[9]~38 (
	.dataa(Mux9),
	.datab(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9~portbdataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[8]~37 ),
	.combout(\dout[9]~38_combout ),
	.cout(\dout[9]~39 ));
defparam \dout[9]~38 .lut_mask = 16'h96DF;
defparam \dout[9]~38 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[10]~40 (
	.dataa(Mux8),
	.datab(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8~portbdataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[9]~39 ),
	.combout(\dout[10]~40_combout ),
	.cout(\dout[10]~41 ));
defparam \dout[10]~40 .lut_mask = 16'h96BF;
defparam \dout[10]~40 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[11]~42 (
	.dataa(Mux7),
	.datab(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7~portbdataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[10]~41 ),
	.combout(\dout[11]~42_combout ),
	.cout(\dout[11]~43 ));
defparam \dout[11]~42 .lut_mask = 16'h96DF;
defparam \dout[11]~42 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[12]~44 (
	.dataa(Mux6),
	.datab(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6~portbdataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[11]~43 ),
	.combout(\dout[12]~44_combout ),
	.cout(\dout[12]~45 ));
defparam \dout[12]~44 .lut_mask = 16'h96BF;
defparam \dout[12]~44 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[13]~46 (
	.dataa(Mux5),
	.datab(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5~portbdataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[12]~45 ),
	.combout(\dout[13]~46_combout ),
	.cout(\dout[13]~47 ));
defparam \dout[13]~46 .lut_mask = 16'h96DF;
defparam \dout[13]~46 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[14]~48 (
	.dataa(Mux4),
	.datab(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4~portbdataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[13]~47 ),
	.combout(\dout[14]~48_combout ),
	.cout(\dout[14]~49 ));
defparam \dout[14]~48 .lut_mask = 16'h96BF;
defparam \dout[14]~48 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[15]~50 (
	.dataa(Mux3),
	.datab(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3~portbdataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[14]~49 ),
	.combout(\dout[15]~50_combout ),
	.cout(\dout[15]~51 ));
defparam \dout[15]~50 .lut_mask = 16'h96DF;
defparam \dout[15]~50 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[16]~52 (
	.dataa(Mux2),
	.datab(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2~portbdataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[15]~51 ),
	.combout(\dout[16]~52_combout ),
	.cout(\dout[16]~53 ));
defparam \dout[16]~52 .lut_mask = 16'h96BF;
defparam \dout[16]~52 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[17]~54 (
	.dataa(Mux1),
	.datab(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1~portbdataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[16]~53 ),
	.combout(\dout[17]~54_combout ),
	.cout(\dout[17]~55 ));
defparam \dout[17]~54 .lut_mask = 16'h96DF;
defparam \dout[17]~54 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[18]~56 (
	.dataa(Mux0),
	.datab(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0~portbdataout ),
	.datac(gnd),
	.datad(gnd),
	.cin(\dout[17]~55 ),
	.combout(\dout[18]~56_combout ),
	.cout());
defparam \dout[18]~56 .lut_mask = 16'h9696;
defparam \dout[18]~56 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout_valid~0 (
	.dataa(reset_n),
	.datab(ena_diff_s_11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\dout_valid~0_combout ),
	.cout());
defparam \dout_valid~0 .lut_mask = 16'hEEEE;
defparam \dout_valid~0 .sum_lutc_input = "datac";

endmodule

module cic_auk_dspip_delay (
	ram_block5a18,
	ram_block5a17,
	ram_block5a16,
	ram_block5a15,
	ram_block5a14,
	ram_block5a13,
	ram_block5a12,
	ram_block5a11,
	ram_block5a10,
	ram_block5a9,
	ram_block5a8,
	ram_block5a7,
	ram_block5a6,
	ram_block5a5,
	ram_block5a4,
	ram_block5a3,
	ram_block5a2,
	ram_block5a1,
	ram_block5a0,
	stall_reg,
	ena_diff_s_1,
	Mux18,
	Mux14,
	Mux13,
	Mux12,
	Mux11,
	Mux10,
	Mux9,
	Mux8,
	Mux7,
	Mux6,
	Mux5,
	Mux4,
	Mux3,
	Mux2,
	Mux1,
	Mux0,
	ena_and_valid,
	Mux17,
	Mux16,
	Mux15,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	ram_block5a18;
output 	ram_block5a17;
output 	ram_block5a16;
output 	ram_block5a15;
output 	ram_block5a14;
output 	ram_block5a13;
output 	ram_block5a12;
output 	ram_block5a11;
output 	ram_block5a10;
output 	ram_block5a9;
output 	ram_block5a8;
output 	ram_block5a7;
output 	ram_block5a6;
output 	ram_block5a5;
output 	ram_block5a4;
output 	ram_block5a3;
output 	ram_block5a2;
output 	ram_block5a1;
output 	ram_block5a0;
input 	stall_reg;
input 	ena_diff_s_1;
input 	Mux18;
input 	Mux14;
input 	Mux13;
input 	Mux12;
input 	Mux11;
input 	Mux10;
input 	Mux9;
input 	Mux8;
input 	Mux7;
input 	Mux6;
input 	Mux5;
input 	Mux4;
input 	Mux3;
input 	Mux2;
input 	Mux1;
input 	Mux0;
input 	ena_and_valid;
input 	Mux17;
input 	Mux16;
input 	Mux15;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0~combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[0]~q ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0~COUT ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1~combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[1]~q ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1~COUT ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~q ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~COUT ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~0_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~0_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~1 ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~2_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~3 ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~4_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~2_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~5 ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[3]~6_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual~combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ;

wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0_PORTBDATAOUT_bus ;

assign ram_block5a18 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18_PORTBDATAOUT_bus [0];

assign ram_block5a17 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17_PORTBDATAOUT_bus [0];

assign ram_block5a16 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16_PORTBDATAOUT_bus [0];

assign ram_block5a15 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15_PORTBDATAOUT_bus [0];

assign ram_block5a14 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14_PORTBDATAOUT_bus [0];

assign ram_block5a13 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13_PORTBDATAOUT_bus [0];

assign ram_block5a12 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12_PORTBDATAOUT_bus [0];

assign ram_block5a11 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11_PORTBDATAOUT_bus [0];

assign ram_block5a10 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10_PORTBDATAOUT_bus [0];

assign ram_block5a9 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9_PORTBDATAOUT_bus [0];

assign ram_block5a8 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8_PORTBDATAOUT_bus [0];

assign ram_block5a7 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7_PORTBDATAOUT_bus [0];

assign ram_block5a6 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6_PORTBDATAOUT_bus [0];

assign ram_block5a5 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5_PORTBDATAOUT_bus [0];

assign ram_block5a4 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4_PORTBDATAOUT_bus [0];

assign ram_block5a3 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3_PORTBDATAOUT_bus [0];

assign ram_block5a2 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2_PORTBDATAOUT_bus [0];

assign ram_block5a1 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1_PORTBDATAOUT_bus [0];

assign ram_block5a0 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0_PORTBDATAOUT_bus [0];

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Mux18}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[0].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_first_bit_number = 18;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_first_bit_number = 18;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Mux17}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[0].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_first_bit_number = 17;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_first_bit_number = 17;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Mux16}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[0].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_first_bit_number = 16;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_first_bit_number = 16;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Mux15}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[0].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_first_bit_number = 15;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_first_bit_number = 15;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Mux14}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[0].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_first_bit_number = 14;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_first_bit_number = 14;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Mux13}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[0].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_first_bit_number = 13;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_first_bit_number = 13;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Mux12}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[0].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_first_bit_number = 12;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_first_bit_number = 12;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Mux11}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[0].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_first_bit_number = 11;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_first_bit_number = 11;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Mux10}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[0].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_first_bit_number = 10;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_first_bit_number = 10;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Mux9}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[0].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_first_bit_number = 9;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_first_bit_number = 9;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Mux8}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[0].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_first_bit_number = 8;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_first_bit_number = 8;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Mux7}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[0].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_first_bit_number = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_first_bit_number = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Mux6}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[0].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_first_bit_number = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_first_bit_number = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Mux5}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[0].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_first_bit_number = 5;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_first_bit_number = 5;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Mux4}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[0].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_first_bit_number = 4;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_first_bit_number = 4;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Mux3}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[0].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_first_bit_number = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_first_bit_number = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Mux2}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[0].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_first_bit_number = 2;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_first_bit_number = 2;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Mux1}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[0].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_first_bit_number = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_first_bit_number = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Mux0}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[0].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_first_bit_number = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_first_bit_number = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .ram_block_type = "auto";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0~combout ),
	.cout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0~COUT ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0 .lut_mask = 16'h55AA;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0 (
	.dataa(stall_reg),
	.datab(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~0_combout ),
	.datac(gnd),
	.datad(ena_diff_s_1),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0 .lut_mask = 16'hFF77;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0_combout ),
	.q(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[0] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0~COUT ),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1~combout ),
	.cout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1~COUT ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1 .lut_mask = 16'h5A5F;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0_combout ),
	.q(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[1] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1~COUT ),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~combout ),
	.cout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~COUT ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2 .lut_mask = 16'h5AAF;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0_combout ),
	.q(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~COUT ),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~0_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~0 .lut_mask = 16'hF0F0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~0 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4 (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena_and_valid),
	.q(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4 .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4 .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~0 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~0_combout ),
	.cout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~1 ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~0 .lut_mask = 16'h55AA;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~2 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~1 ),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~2_combout ),
	.cout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~3 ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~2 .lut_mask = 16'h5A5F;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1 .lut_mask = 16'hAAFF;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena_and_valid),
	.q(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~4 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~3 ),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~4_combout ),
	.cout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~5 ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~4 .lut_mask = 16'h5AAF;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~2 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~2_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~2 .lut_mask = 16'hAAFF;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~2 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena_and_valid),
	.q(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[3]~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~5 ),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[3]~6_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[3]~6 .lut_mask = 16'hF0F0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[3]~6 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[3]~6_combout ),
	.datab(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datac(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datad(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual .lut_mask = 16'hFEFF;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0 .lut_mask = 16'hAAFF;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena_and_valid),
	.q(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .power_up = "low";

endmodule

module cic_auk_dspip_differentiator_1 (
	dout_0,
	dout_1,
	dout_2,
	dout_3,
	dout_4,
	dout_5,
	dout_6,
	dout_7,
	dout_8,
	dout_9,
	dout_10,
	dout_11,
	dout_12,
	dout_13,
	dout_14,
	dout_15,
	dout_16,
	dout_17,
	dout_18,
	dout_01,
	dout_19,
	dout_21,
	dout_31,
	dout_41,
	dout_51,
	dout_61,
	dout_71,
	dout_81,
	dout_91,
	dout_101,
	dout_111,
	dout_121,
	dout_131,
	dout_141,
	dout_151,
	dout_161,
	dout_171,
	dout_181,
	stall_reg,
	dout_valid1,
	ena_diff_s_1,
	dout_valid2,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dout_0;
output 	dout_1;
output 	dout_2;
output 	dout_3;
output 	dout_4;
output 	dout_5;
output 	dout_6;
output 	dout_7;
output 	dout_8;
output 	dout_9;
output 	dout_10;
output 	dout_11;
output 	dout_12;
output 	dout_13;
output 	dout_14;
output 	dout_15;
output 	dout_16;
output 	dout_17;
output 	dout_18;
input 	dout_01;
input 	dout_19;
input 	dout_21;
input 	dout_31;
input 	dout_41;
input 	dout_51;
input 	dout_61;
input 	dout_71;
input 	dout_81;
input 	dout_91;
input 	dout_101;
input 	dout_111;
input 	dout_121;
input 	dout_131;
input 	dout_141;
input 	dout_151;
input 	dout_161;
input 	dout_171;
input 	dout_181;
input 	stall_reg;
output 	dout_valid1;
input 	ena_diff_s_1;
input 	dout_valid2;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0~portbdataout ;
wire \ena_and_valid~combout ;
wire \dout[0]~19_combout ;
wire \dout[1]~21_combout ;
wire \dout[0]~20 ;
wire \dout[1]~22_combout ;
wire \dout[1]~23 ;
wire \dout[2]~24_combout ;
wire \dout[2]~25 ;
wire \dout[3]~26_combout ;
wire \dout[3]~27 ;
wire \dout[4]~28_combout ;
wire \dout[4]~29 ;
wire \dout[5]~30_combout ;
wire \dout[5]~31 ;
wire \dout[6]~32_combout ;
wire \dout[6]~33 ;
wire \dout[7]~34_combout ;
wire \dout[7]~35 ;
wire \dout[8]~36_combout ;
wire \dout[8]~37 ;
wire \dout[9]~38_combout ;
wire \dout[9]~39 ;
wire \dout[10]~40_combout ;
wire \dout[10]~41 ;
wire \dout[11]~42_combout ;
wire \dout[11]~43 ;
wire \dout[12]~44_combout ;
wire \dout[12]~45 ;
wire \dout[13]~46_combout ;
wire \dout[13]~47 ;
wire \dout[14]~48_combout ;
wire \dout[14]~49 ;
wire \dout[15]~50_combout ;
wire \dout[15]~51 ;
wire \dout[16]~52_combout ;
wire \dout[16]~53 ;
wire \dout[17]~54_combout ;
wire \dout[17]~55 ;
wire \dout[18]~56_combout ;
wire \dout_valid~0_combout ;


cic_auk_dspip_delay_1 \glogic:u0 (
	.ram_block5a18(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18~portbdataout ),
	.dout_0(dout_01),
	.ram_block5a17(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17~portbdataout ),
	.dout_1(dout_19),
	.ram_block5a16(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16~portbdataout ),
	.dout_2(dout_21),
	.ram_block5a15(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15~portbdataout ),
	.dout_3(dout_31),
	.ram_block5a14(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14~portbdataout ),
	.dout_4(dout_41),
	.ram_block5a13(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13~portbdataout ),
	.dout_5(dout_51),
	.ram_block5a12(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12~portbdataout ),
	.dout_6(dout_61),
	.ram_block5a11(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11~portbdataout ),
	.dout_7(dout_71),
	.ram_block5a10(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10~portbdataout ),
	.dout_8(dout_81),
	.ram_block5a9(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9~portbdataout ),
	.dout_9(dout_91),
	.ram_block5a8(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8~portbdataout ),
	.dout_10(dout_101),
	.ram_block5a7(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7~portbdataout ),
	.dout_11(dout_111),
	.ram_block5a6(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6~portbdataout ),
	.dout_12(dout_121),
	.ram_block5a5(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5~portbdataout ),
	.dout_13(dout_131),
	.ram_block5a4(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4~portbdataout ),
	.dout_14(dout_141),
	.ram_block5a3(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3~portbdataout ),
	.dout_15(dout_151),
	.ram_block5a2(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2~portbdataout ),
	.dout_16(dout_161),
	.ram_block5a1(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1~portbdataout ),
	.dout_17(dout_171),
	.ram_block5a0(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0~portbdataout ),
	.dout_18(dout_181),
	.stall_reg(stall_reg),
	.dout_valid(dout_valid2),
	.ena_and_valid(\ena_and_valid~combout ),
	.clk(clk),
	.reset_n(reset_n));

fiftyfivenm_lcell_comb ena_and_valid(
	.dataa(stall_reg),
	.datab(gnd),
	.datac(gnd),
	.datad(dout_valid2),
	.cin(gnd),
	.combout(\ena_and_valid~combout ),
	.cout());
defparam ena_and_valid.lut_mask = 16'hFF55;
defparam ena_and_valid.sum_lutc_input = "datac";

dffeas \dout[0] (
	.clk(clk),
	.d(\dout[0]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[1]~21_combout ),
	.q(dout_0),
	.prn(vcc));
defparam \dout[0] .is_wysiwyg = "true";
defparam \dout[0] .power_up = "low";

dffeas \dout[1] (
	.clk(clk),
	.d(\dout[1]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[1]~21_combout ),
	.q(dout_1),
	.prn(vcc));
defparam \dout[1] .is_wysiwyg = "true";
defparam \dout[1] .power_up = "low";

dffeas \dout[2] (
	.clk(clk),
	.d(\dout[2]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[1]~21_combout ),
	.q(dout_2),
	.prn(vcc));
defparam \dout[2] .is_wysiwyg = "true";
defparam \dout[2] .power_up = "low";

dffeas \dout[3] (
	.clk(clk),
	.d(\dout[3]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[1]~21_combout ),
	.q(dout_3),
	.prn(vcc));
defparam \dout[3] .is_wysiwyg = "true";
defparam \dout[3] .power_up = "low";

dffeas \dout[4] (
	.clk(clk),
	.d(\dout[4]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[1]~21_combout ),
	.q(dout_4),
	.prn(vcc));
defparam \dout[4] .is_wysiwyg = "true";
defparam \dout[4] .power_up = "low";

dffeas \dout[5] (
	.clk(clk),
	.d(\dout[5]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[1]~21_combout ),
	.q(dout_5),
	.prn(vcc));
defparam \dout[5] .is_wysiwyg = "true";
defparam \dout[5] .power_up = "low";

dffeas \dout[6] (
	.clk(clk),
	.d(\dout[6]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[1]~21_combout ),
	.q(dout_6),
	.prn(vcc));
defparam \dout[6] .is_wysiwyg = "true";
defparam \dout[6] .power_up = "low";

dffeas \dout[7] (
	.clk(clk),
	.d(\dout[7]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[1]~21_combout ),
	.q(dout_7),
	.prn(vcc));
defparam \dout[7] .is_wysiwyg = "true";
defparam \dout[7] .power_up = "low";

dffeas \dout[8] (
	.clk(clk),
	.d(\dout[8]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[1]~21_combout ),
	.q(dout_8),
	.prn(vcc));
defparam \dout[8] .is_wysiwyg = "true";
defparam \dout[8] .power_up = "low";

dffeas \dout[9] (
	.clk(clk),
	.d(\dout[9]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[1]~21_combout ),
	.q(dout_9),
	.prn(vcc));
defparam \dout[9] .is_wysiwyg = "true";
defparam \dout[9] .power_up = "low";

dffeas \dout[10] (
	.clk(clk),
	.d(\dout[10]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[1]~21_combout ),
	.q(dout_10),
	.prn(vcc));
defparam \dout[10] .is_wysiwyg = "true";
defparam \dout[10] .power_up = "low";

dffeas \dout[11] (
	.clk(clk),
	.d(\dout[11]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[1]~21_combout ),
	.q(dout_11),
	.prn(vcc));
defparam \dout[11] .is_wysiwyg = "true";
defparam \dout[11] .power_up = "low";

dffeas \dout[12] (
	.clk(clk),
	.d(\dout[12]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[1]~21_combout ),
	.q(dout_12),
	.prn(vcc));
defparam \dout[12] .is_wysiwyg = "true";
defparam \dout[12] .power_up = "low";

dffeas \dout[13] (
	.clk(clk),
	.d(\dout[13]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[1]~21_combout ),
	.q(dout_13),
	.prn(vcc));
defparam \dout[13] .is_wysiwyg = "true";
defparam \dout[13] .power_up = "low";

dffeas \dout[14] (
	.clk(clk),
	.d(\dout[14]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[1]~21_combout ),
	.q(dout_14),
	.prn(vcc));
defparam \dout[14] .is_wysiwyg = "true";
defparam \dout[14] .power_up = "low";

dffeas \dout[15] (
	.clk(clk),
	.d(\dout[15]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[1]~21_combout ),
	.q(dout_15),
	.prn(vcc));
defparam \dout[15] .is_wysiwyg = "true";
defparam \dout[15] .power_up = "low";

dffeas \dout[16] (
	.clk(clk),
	.d(\dout[16]~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[1]~21_combout ),
	.q(dout_16),
	.prn(vcc));
defparam \dout[16] .is_wysiwyg = "true";
defparam \dout[16] .power_up = "low";

dffeas \dout[17] (
	.clk(clk),
	.d(\dout[17]~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[1]~21_combout ),
	.q(dout_17),
	.prn(vcc));
defparam \dout[17] .is_wysiwyg = "true";
defparam \dout[17] .power_up = "low";

dffeas \dout[18] (
	.clk(clk),
	.d(\dout[18]~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[1]~21_combout ),
	.q(dout_18),
	.prn(vcc));
defparam \dout[18] .is_wysiwyg = "true";
defparam \dout[18] .power_up = "low";

dffeas dout_valid(
	.clk(clk),
	.d(\dout_valid~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena_diff_s_1),
	.q(dout_valid1),
	.prn(vcc));
defparam dout_valid.is_wysiwyg = "true";
defparam dout_valid.power_up = "low";

fiftyfivenm_lcell_comb \dout[0]~19 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18~portbdataout ),
	.datab(dout_01),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\dout[0]~19_combout ),
	.cout(\dout[0]~20 ));
defparam \dout[0]~19 .lut_mask = 16'h66DD;
defparam \dout[0]~19 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dout[1]~21 (
	.dataa(reset_n),
	.datab(stall_reg),
	.datac(gnd),
	.datad(dout_valid2),
	.cin(gnd),
	.combout(\dout[1]~21_combout ),
	.cout());
defparam \dout[1]~21 .lut_mask = 16'hFF77;
defparam \dout[1]~21 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dout[1]~22 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17~portbdataout ),
	.datab(dout_19),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[0]~20 ),
	.combout(\dout[1]~22_combout ),
	.cout(\dout[1]~23 ));
defparam \dout[1]~22 .lut_mask = 16'h96BF;
defparam \dout[1]~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[2]~24 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16~portbdataout ),
	.datab(dout_21),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[1]~23 ),
	.combout(\dout[2]~24_combout ),
	.cout(\dout[2]~25 ));
defparam \dout[2]~24 .lut_mask = 16'h96DF;
defparam \dout[2]~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[3]~26 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15~portbdataout ),
	.datab(dout_31),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[2]~25 ),
	.combout(\dout[3]~26_combout ),
	.cout(\dout[3]~27 ));
defparam \dout[3]~26 .lut_mask = 16'h96BF;
defparam \dout[3]~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[4]~28 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14~portbdataout ),
	.datab(dout_41),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[3]~27 ),
	.combout(\dout[4]~28_combout ),
	.cout(\dout[4]~29 ));
defparam \dout[4]~28 .lut_mask = 16'h96DF;
defparam \dout[4]~28 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[5]~30 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13~portbdataout ),
	.datab(dout_51),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[4]~29 ),
	.combout(\dout[5]~30_combout ),
	.cout(\dout[5]~31 ));
defparam \dout[5]~30 .lut_mask = 16'h96BF;
defparam \dout[5]~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[6]~32 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12~portbdataout ),
	.datab(dout_61),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[5]~31 ),
	.combout(\dout[6]~32_combout ),
	.cout(\dout[6]~33 ));
defparam \dout[6]~32 .lut_mask = 16'h96DF;
defparam \dout[6]~32 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[7]~34 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11~portbdataout ),
	.datab(dout_71),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[6]~33 ),
	.combout(\dout[7]~34_combout ),
	.cout(\dout[7]~35 ));
defparam \dout[7]~34 .lut_mask = 16'h96BF;
defparam \dout[7]~34 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[8]~36 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10~portbdataout ),
	.datab(dout_81),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[7]~35 ),
	.combout(\dout[8]~36_combout ),
	.cout(\dout[8]~37 ));
defparam \dout[8]~36 .lut_mask = 16'h96DF;
defparam \dout[8]~36 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[9]~38 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9~portbdataout ),
	.datab(dout_91),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[8]~37 ),
	.combout(\dout[9]~38_combout ),
	.cout(\dout[9]~39 ));
defparam \dout[9]~38 .lut_mask = 16'h96BF;
defparam \dout[9]~38 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[10]~40 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8~portbdataout ),
	.datab(dout_101),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[9]~39 ),
	.combout(\dout[10]~40_combout ),
	.cout(\dout[10]~41 ));
defparam \dout[10]~40 .lut_mask = 16'h96DF;
defparam \dout[10]~40 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[11]~42 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7~portbdataout ),
	.datab(dout_111),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[10]~41 ),
	.combout(\dout[11]~42_combout ),
	.cout(\dout[11]~43 ));
defparam \dout[11]~42 .lut_mask = 16'h96BF;
defparam \dout[11]~42 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[12]~44 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6~portbdataout ),
	.datab(dout_121),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[11]~43 ),
	.combout(\dout[12]~44_combout ),
	.cout(\dout[12]~45 ));
defparam \dout[12]~44 .lut_mask = 16'h96DF;
defparam \dout[12]~44 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[13]~46 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5~portbdataout ),
	.datab(dout_131),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[12]~45 ),
	.combout(\dout[13]~46_combout ),
	.cout(\dout[13]~47 ));
defparam \dout[13]~46 .lut_mask = 16'h96BF;
defparam \dout[13]~46 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[14]~48 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4~portbdataout ),
	.datab(dout_141),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[13]~47 ),
	.combout(\dout[14]~48_combout ),
	.cout(\dout[14]~49 ));
defparam \dout[14]~48 .lut_mask = 16'h96DF;
defparam \dout[14]~48 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[15]~50 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3~portbdataout ),
	.datab(dout_151),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[14]~49 ),
	.combout(\dout[15]~50_combout ),
	.cout(\dout[15]~51 ));
defparam \dout[15]~50 .lut_mask = 16'h96BF;
defparam \dout[15]~50 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[16]~52 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2~portbdataout ),
	.datab(dout_161),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[15]~51 ),
	.combout(\dout[16]~52_combout ),
	.cout(\dout[16]~53 ));
defparam \dout[16]~52 .lut_mask = 16'h96DF;
defparam \dout[16]~52 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[17]~54 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1~portbdataout ),
	.datab(dout_171),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[16]~53 ),
	.combout(\dout[17]~54_combout ),
	.cout(\dout[17]~55 ));
defparam \dout[17]~54 .lut_mask = 16'h96BF;
defparam \dout[17]~54 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[18]~56 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0~portbdataout ),
	.datab(dout_181),
	.datac(gnd),
	.datad(gnd),
	.cin(\dout[17]~55 ),
	.combout(\dout[18]~56_combout ),
	.cout());
defparam \dout[18]~56 .lut_mask = 16'h9696;
defparam \dout[18]~56 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout_valid~0 (
	.dataa(reset_n),
	.datab(dout_valid2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\dout_valid~0_combout ),
	.cout());
defparam \dout_valid~0 .lut_mask = 16'hEEEE;
defparam \dout_valid~0 .sum_lutc_input = "datac";

endmodule

module cic_auk_dspip_delay_1 (
	ram_block5a18,
	dout_0,
	ram_block5a17,
	dout_1,
	ram_block5a16,
	dout_2,
	ram_block5a15,
	dout_3,
	ram_block5a14,
	dout_4,
	ram_block5a13,
	dout_5,
	ram_block5a12,
	dout_6,
	ram_block5a11,
	dout_7,
	ram_block5a10,
	dout_8,
	ram_block5a9,
	dout_9,
	ram_block5a8,
	dout_10,
	ram_block5a7,
	dout_11,
	ram_block5a6,
	dout_12,
	ram_block5a5,
	dout_13,
	ram_block5a4,
	dout_14,
	ram_block5a3,
	dout_15,
	ram_block5a2,
	dout_16,
	ram_block5a1,
	dout_17,
	ram_block5a0,
	dout_18,
	stall_reg,
	dout_valid,
	ena_and_valid,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	ram_block5a18;
input 	dout_0;
output 	ram_block5a17;
input 	dout_1;
output 	ram_block5a16;
input 	dout_2;
output 	ram_block5a15;
input 	dout_3;
output 	ram_block5a14;
input 	dout_4;
output 	ram_block5a13;
input 	dout_5;
output 	ram_block5a12;
input 	dout_6;
output 	ram_block5a11;
input 	dout_7;
output 	ram_block5a10;
input 	dout_8;
output 	ram_block5a9;
input 	dout_9;
output 	ram_block5a8;
input 	dout_10;
output 	ram_block5a7;
input 	dout_11;
output 	ram_block5a6;
input 	dout_12;
output 	ram_block5a5;
input 	dout_13;
output 	ram_block5a4;
input 	dout_14;
output 	ram_block5a3;
input 	dout_15;
output 	ram_block5a2;
input 	dout_16;
output 	ram_block5a1;
input 	dout_17;
output 	ram_block5a0;
input 	dout_18;
input 	stall_reg;
input 	dout_valid;
input 	ena_and_valid;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0~combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[0]~q ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0~COUT ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1~combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[1]~q ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1~COUT ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~q ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~COUT ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~0_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~0_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~1 ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~2_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~3 ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~4_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~2_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~5 ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[3]~6_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual~combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ;

wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0_PORTBDATAOUT_bus ;

assign ram_block5a18 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18_PORTBDATAOUT_bus [0];

assign ram_block5a17 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17_PORTBDATAOUT_bus [0];

assign ram_block5a16 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16_PORTBDATAOUT_bus [0];

assign ram_block5a15 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15_PORTBDATAOUT_bus [0];

assign ram_block5a14 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14_PORTBDATAOUT_bus [0];

assign ram_block5a13 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13_PORTBDATAOUT_bus [0];

assign ram_block5a12 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12_PORTBDATAOUT_bus [0];

assign ram_block5a11 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11_PORTBDATAOUT_bus [0];

assign ram_block5a10 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10_PORTBDATAOUT_bus [0];

assign ram_block5a9 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9_PORTBDATAOUT_bus [0];

assign ram_block5a8 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8_PORTBDATAOUT_bus [0];

assign ram_block5a7 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7_PORTBDATAOUT_bus [0];

assign ram_block5a6 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6_PORTBDATAOUT_bus [0];

assign ram_block5a5 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5_PORTBDATAOUT_bus [0];

assign ram_block5a4 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4_PORTBDATAOUT_bus [0];

assign ram_block5a3 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3_PORTBDATAOUT_bus [0];

assign ram_block5a2 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2_PORTBDATAOUT_bus [0];

assign ram_block5a1 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1_PORTBDATAOUT_bus [0];

assign ram_block5a0 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0_PORTBDATAOUT_bus [0];

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_0}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[1].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_first_bit_number = 18;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_first_bit_number = 18;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_1}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[1].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_first_bit_number = 17;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_first_bit_number = 17;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_2}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[1].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_first_bit_number = 16;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_first_bit_number = 16;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_3}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[1].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_first_bit_number = 15;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_first_bit_number = 15;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_4}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[1].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_first_bit_number = 14;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_first_bit_number = 14;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_5}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[1].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_first_bit_number = 13;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_first_bit_number = 13;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_6}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[1].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_first_bit_number = 12;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_first_bit_number = 12;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_7}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[1].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_first_bit_number = 11;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_first_bit_number = 11;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_8}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[1].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_first_bit_number = 10;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_first_bit_number = 10;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_9}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[1].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_first_bit_number = 9;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_first_bit_number = 9;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_10}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[1].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_first_bit_number = 8;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_first_bit_number = 8;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_11}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[1].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_first_bit_number = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_first_bit_number = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_12}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[1].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_first_bit_number = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_first_bit_number = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_13}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[1].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_first_bit_number = 5;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_first_bit_number = 5;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_14}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[1].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_first_bit_number = 4;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_first_bit_number = 4;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_15}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[1].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_first_bit_number = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_first_bit_number = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_16}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[1].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_first_bit_number = 2;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_first_bit_number = 2;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_17}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[1].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_first_bit_number = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_first_bit_number = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_18}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[1].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_first_bit_number = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_first_bit_number = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .ram_block_type = "auto";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0~combout ),
	.cout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0~COUT ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0 .lut_mask = 16'h55AA;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0 (
	.dataa(stall_reg),
	.datab(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~0_combout ),
	.datac(gnd),
	.datad(dout_valid),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0 .lut_mask = 16'hFF77;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0_combout ),
	.q(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[0] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0~COUT ),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1~combout ),
	.cout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1~COUT ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1 .lut_mask = 16'h5A5F;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0_combout ),
	.q(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[1] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1~COUT ),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~combout ),
	.cout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~COUT ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2 .lut_mask = 16'h5AAF;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0_combout ),
	.q(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~COUT ),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~0_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~0 .lut_mask = 16'hF0F0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~0 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4 (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena_and_valid),
	.q(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4 .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4 .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~0 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~0_combout ),
	.cout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~1 ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~0 .lut_mask = 16'h55AA;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~2 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~1 ),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~2_combout ),
	.cout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~3 ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~2 .lut_mask = 16'h5A5F;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1 .lut_mask = 16'hAAFF;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena_and_valid),
	.q(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~4 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~3 ),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~4_combout ),
	.cout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~5 ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~4 .lut_mask = 16'h5AAF;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~2 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~2_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~2 .lut_mask = 16'hAAFF;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~2 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena_and_valid),
	.q(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[3]~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~5 ),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[3]~6_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[3]~6 .lut_mask = 16'hF0F0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[3]~6 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[3]~6_combout ),
	.datab(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datac(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datad(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual .lut_mask = 16'hFEFF;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0 .lut_mask = 16'hAAFF;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena_and_valid),
	.q(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .power_up = "low";

endmodule

module cic_auk_dspip_differentiator_2 (
	dout_0,
	dout_1,
	dout_2,
	dout_3,
	dout_4,
	dout_5,
	dout_6,
	dout_7,
	dout_8,
	dout_9,
	dout_10,
	dout_11,
	dout_12,
	dout_13,
	dout_14,
	dout_15,
	dout_16,
	dout_17,
	dout_18,
	dout_01,
	dout_19,
	dout_21,
	dout_31,
	dout_41,
	dout_51,
	dout_61,
	dout_71,
	dout_81,
	dout_91,
	dout_101,
	dout_111,
	dout_121,
	dout_131,
	dout_141,
	dout_151,
	dout_161,
	dout_171,
	dout_181,
	stall_reg,
	dout_valid1,
	dout_valid2,
	ena_diff_s_1,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dout_0;
output 	dout_1;
output 	dout_2;
output 	dout_3;
output 	dout_4;
output 	dout_5;
output 	dout_6;
output 	dout_7;
output 	dout_8;
output 	dout_9;
output 	dout_10;
output 	dout_11;
output 	dout_12;
output 	dout_13;
output 	dout_14;
output 	dout_15;
output 	dout_16;
output 	dout_17;
output 	dout_18;
input 	dout_01;
input 	dout_19;
input 	dout_21;
input 	dout_31;
input 	dout_41;
input 	dout_51;
input 	dout_61;
input 	dout_71;
input 	dout_81;
input 	dout_91;
input 	dout_101;
input 	dout_111;
input 	dout_121;
input 	dout_131;
input 	dout_141;
input 	dout_151;
input 	dout_161;
input 	dout_171;
input 	dout_181;
input 	stall_reg;
output 	dout_valid1;
input 	dout_valid2;
input 	ena_diff_s_1;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1~portbdataout ;
wire \glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0~portbdataout ;
wire \ena_and_valid~combout ;
wire \dout[0]~19_combout ;
wire \dout[3]~21_combout ;
wire \dout[0]~20 ;
wire \dout[1]~22_combout ;
wire \dout[1]~23 ;
wire \dout[2]~24_combout ;
wire \dout[2]~25 ;
wire \dout[3]~26_combout ;
wire \dout[3]~27 ;
wire \dout[4]~28_combout ;
wire \dout[4]~29 ;
wire \dout[5]~30_combout ;
wire \dout[5]~31 ;
wire \dout[6]~32_combout ;
wire \dout[6]~33 ;
wire \dout[7]~34_combout ;
wire \dout[7]~35 ;
wire \dout[8]~36_combout ;
wire \dout[8]~37 ;
wire \dout[9]~38_combout ;
wire \dout[9]~39 ;
wire \dout[10]~40_combout ;
wire \dout[10]~41 ;
wire \dout[11]~42_combout ;
wire \dout[11]~43 ;
wire \dout[12]~44_combout ;
wire \dout[12]~45 ;
wire \dout[13]~46_combout ;
wire \dout[13]~47 ;
wire \dout[14]~48_combout ;
wire \dout[14]~49 ;
wire \dout[15]~50_combout ;
wire \dout[15]~51 ;
wire \dout[16]~52_combout ;
wire \dout[16]~53 ;
wire \dout[17]~54_combout ;
wire \dout[17]~55 ;
wire \dout[18]~56_combout ;
wire \dout_valid~0_combout ;


cic_auk_dspip_delay_2 \glogic:u0 (
	.ram_block5a18(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18~portbdataout ),
	.dout_0(dout_01),
	.ram_block5a17(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17~portbdataout ),
	.dout_1(dout_19),
	.ram_block5a16(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16~portbdataout ),
	.dout_2(dout_21),
	.ram_block5a15(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15~portbdataout ),
	.dout_3(dout_31),
	.ram_block5a14(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14~portbdataout ),
	.dout_4(dout_41),
	.ram_block5a13(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13~portbdataout ),
	.dout_5(dout_51),
	.ram_block5a12(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12~portbdataout ),
	.dout_6(dout_61),
	.ram_block5a11(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11~portbdataout ),
	.dout_7(dout_71),
	.ram_block5a10(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10~portbdataout ),
	.dout_8(dout_81),
	.ram_block5a9(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9~portbdataout ),
	.dout_9(dout_91),
	.ram_block5a8(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8~portbdataout ),
	.dout_10(dout_101),
	.ram_block5a7(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7~portbdataout ),
	.dout_11(dout_111),
	.ram_block5a6(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6~portbdataout ),
	.dout_12(dout_121),
	.ram_block5a5(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5~portbdataout ),
	.dout_13(dout_131),
	.ram_block5a4(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4~portbdataout ),
	.dout_14(dout_141),
	.ram_block5a3(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3~portbdataout ),
	.dout_15(dout_151),
	.ram_block5a2(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2~portbdataout ),
	.dout_16(dout_161),
	.ram_block5a1(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1~portbdataout ),
	.dout_17(dout_171),
	.ram_block5a0(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0~portbdataout ),
	.dout_18(dout_181),
	.stall_reg(stall_reg),
	.dout_valid(dout_valid2),
	.ena_and_valid(\ena_and_valid~combout ),
	.clk(clk),
	.reset_n(reset_n));

fiftyfivenm_lcell_comb ena_and_valid(
	.dataa(stall_reg),
	.datab(gnd),
	.datac(gnd),
	.datad(dout_valid2),
	.cin(gnd),
	.combout(\ena_and_valid~combout ),
	.cout());
defparam ena_and_valid.lut_mask = 16'hFF55;
defparam ena_and_valid.sum_lutc_input = "datac";

dffeas \dout[0] (
	.clk(clk),
	.d(\dout[0]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[3]~21_combout ),
	.q(dout_0),
	.prn(vcc));
defparam \dout[0] .is_wysiwyg = "true";
defparam \dout[0] .power_up = "low";

dffeas \dout[1] (
	.clk(clk),
	.d(\dout[1]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[3]~21_combout ),
	.q(dout_1),
	.prn(vcc));
defparam \dout[1] .is_wysiwyg = "true";
defparam \dout[1] .power_up = "low";

dffeas \dout[2] (
	.clk(clk),
	.d(\dout[2]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[3]~21_combout ),
	.q(dout_2),
	.prn(vcc));
defparam \dout[2] .is_wysiwyg = "true";
defparam \dout[2] .power_up = "low";

dffeas \dout[3] (
	.clk(clk),
	.d(\dout[3]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[3]~21_combout ),
	.q(dout_3),
	.prn(vcc));
defparam \dout[3] .is_wysiwyg = "true";
defparam \dout[3] .power_up = "low";

dffeas \dout[4] (
	.clk(clk),
	.d(\dout[4]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[3]~21_combout ),
	.q(dout_4),
	.prn(vcc));
defparam \dout[4] .is_wysiwyg = "true";
defparam \dout[4] .power_up = "low";

dffeas \dout[5] (
	.clk(clk),
	.d(\dout[5]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[3]~21_combout ),
	.q(dout_5),
	.prn(vcc));
defparam \dout[5] .is_wysiwyg = "true";
defparam \dout[5] .power_up = "low";

dffeas \dout[6] (
	.clk(clk),
	.d(\dout[6]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[3]~21_combout ),
	.q(dout_6),
	.prn(vcc));
defparam \dout[6] .is_wysiwyg = "true";
defparam \dout[6] .power_up = "low";

dffeas \dout[7] (
	.clk(clk),
	.d(\dout[7]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[3]~21_combout ),
	.q(dout_7),
	.prn(vcc));
defparam \dout[7] .is_wysiwyg = "true";
defparam \dout[7] .power_up = "low";

dffeas \dout[8] (
	.clk(clk),
	.d(\dout[8]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[3]~21_combout ),
	.q(dout_8),
	.prn(vcc));
defparam \dout[8] .is_wysiwyg = "true";
defparam \dout[8] .power_up = "low";

dffeas \dout[9] (
	.clk(clk),
	.d(\dout[9]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[3]~21_combout ),
	.q(dout_9),
	.prn(vcc));
defparam \dout[9] .is_wysiwyg = "true";
defparam \dout[9] .power_up = "low";

dffeas \dout[10] (
	.clk(clk),
	.d(\dout[10]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[3]~21_combout ),
	.q(dout_10),
	.prn(vcc));
defparam \dout[10] .is_wysiwyg = "true";
defparam \dout[10] .power_up = "low";

dffeas \dout[11] (
	.clk(clk),
	.d(\dout[11]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[3]~21_combout ),
	.q(dout_11),
	.prn(vcc));
defparam \dout[11] .is_wysiwyg = "true";
defparam \dout[11] .power_up = "low";

dffeas \dout[12] (
	.clk(clk),
	.d(\dout[12]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[3]~21_combout ),
	.q(dout_12),
	.prn(vcc));
defparam \dout[12] .is_wysiwyg = "true";
defparam \dout[12] .power_up = "low";

dffeas \dout[13] (
	.clk(clk),
	.d(\dout[13]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[3]~21_combout ),
	.q(dout_13),
	.prn(vcc));
defparam \dout[13] .is_wysiwyg = "true";
defparam \dout[13] .power_up = "low";

dffeas \dout[14] (
	.clk(clk),
	.d(\dout[14]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[3]~21_combout ),
	.q(dout_14),
	.prn(vcc));
defparam \dout[14] .is_wysiwyg = "true";
defparam \dout[14] .power_up = "low";

dffeas \dout[15] (
	.clk(clk),
	.d(\dout[15]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[3]~21_combout ),
	.q(dout_15),
	.prn(vcc));
defparam \dout[15] .is_wysiwyg = "true";
defparam \dout[15] .power_up = "low";

dffeas \dout[16] (
	.clk(clk),
	.d(\dout[16]~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[3]~21_combout ),
	.q(dout_16),
	.prn(vcc));
defparam \dout[16] .is_wysiwyg = "true";
defparam \dout[16] .power_up = "low";

dffeas \dout[17] (
	.clk(clk),
	.d(\dout[17]~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[3]~21_combout ),
	.q(dout_17),
	.prn(vcc));
defparam \dout[17] .is_wysiwyg = "true";
defparam \dout[17] .power_up = "low";

dffeas \dout[18] (
	.clk(clk),
	.d(\dout[18]~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\dout[3]~21_combout ),
	.q(dout_18),
	.prn(vcc));
defparam \dout[18] .is_wysiwyg = "true";
defparam \dout[18] .power_up = "low";

dffeas dout_valid(
	.clk(clk),
	.d(\dout_valid~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena_diff_s_1),
	.q(dout_valid1),
	.prn(vcc));
defparam dout_valid.is_wysiwyg = "true";
defparam dout_valid.power_up = "low";

fiftyfivenm_lcell_comb \dout[0]~19 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18~portbdataout ),
	.datab(dout_01),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\dout[0]~19_combout ),
	.cout(\dout[0]~20 ));
defparam \dout[0]~19 .lut_mask = 16'h66DD;
defparam \dout[0]~19 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dout[3]~21 (
	.dataa(reset_n),
	.datab(stall_reg),
	.datac(gnd),
	.datad(dout_valid2),
	.cin(gnd),
	.combout(\dout[3]~21_combout ),
	.cout());
defparam \dout[3]~21 .lut_mask = 16'hFF77;
defparam \dout[3]~21 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dout[1]~22 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17~portbdataout ),
	.datab(dout_19),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[0]~20 ),
	.combout(\dout[1]~22_combout ),
	.cout(\dout[1]~23 ));
defparam \dout[1]~22 .lut_mask = 16'h96BF;
defparam \dout[1]~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[2]~24 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16~portbdataout ),
	.datab(dout_21),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[1]~23 ),
	.combout(\dout[2]~24_combout ),
	.cout(\dout[2]~25 ));
defparam \dout[2]~24 .lut_mask = 16'h96DF;
defparam \dout[2]~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[3]~26 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15~portbdataout ),
	.datab(dout_31),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[2]~25 ),
	.combout(\dout[3]~26_combout ),
	.cout(\dout[3]~27 ));
defparam \dout[3]~26 .lut_mask = 16'h96BF;
defparam \dout[3]~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[4]~28 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14~portbdataout ),
	.datab(dout_41),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[3]~27 ),
	.combout(\dout[4]~28_combout ),
	.cout(\dout[4]~29 ));
defparam \dout[4]~28 .lut_mask = 16'h96DF;
defparam \dout[4]~28 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[5]~30 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13~portbdataout ),
	.datab(dout_51),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[4]~29 ),
	.combout(\dout[5]~30_combout ),
	.cout(\dout[5]~31 ));
defparam \dout[5]~30 .lut_mask = 16'h96BF;
defparam \dout[5]~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[6]~32 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12~portbdataout ),
	.datab(dout_61),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[5]~31 ),
	.combout(\dout[6]~32_combout ),
	.cout(\dout[6]~33 ));
defparam \dout[6]~32 .lut_mask = 16'h96DF;
defparam \dout[6]~32 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[7]~34 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11~portbdataout ),
	.datab(dout_71),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[6]~33 ),
	.combout(\dout[7]~34_combout ),
	.cout(\dout[7]~35 ));
defparam \dout[7]~34 .lut_mask = 16'h96BF;
defparam \dout[7]~34 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[8]~36 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10~portbdataout ),
	.datab(dout_81),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[7]~35 ),
	.combout(\dout[8]~36_combout ),
	.cout(\dout[8]~37 ));
defparam \dout[8]~36 .lut_mask = 16'h96DF;
defparam \dout[8]~36 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[9]~38 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9~portbdataout ),
	.datab(dout_91),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[8]~37 ),
	.combout(\dout[9]~38_combout ),
	.cout(\dout[9]~39 ));
defparam \dout[9]~38 .lut_mask = 16'h96BF;
defparam \dout[9]~38 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[10]~40 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8~portbdataout ),
	.datab(dout_101),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[9]~39 ),
	.combout(\dout[10]~40_combout ),
	.cout(\dout[10]~41 ));
defparam \dout[10]~40 .lut_mask = 16'h96DF;
defparam \dout[10]~40 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[11]~42 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7~portbdataout ),
	.datab(dout_111),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[10]~41 ),
	.combout(\dout[11]~42_combout ),
	.cout(\dout[11]~43 ));
defparam \dout[11]~42 .lut_mask = 16'h96BF;
defparam \dout[11]~42 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[12]~44 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6~portbdataout ),
	.datab(dout_121),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[11]~43 ),
	.combout(\dout[12]~44_combout ),
	.cout(\dout[12]~45 ));
defparam \dout[12]~44 .lut_mask = 16'h96DF;
defparam \dout[12]~44 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[13]~46 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5~portbdataout ),
	.datab(dout_131),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[12]~45 ),
	.combout(\dout[13]~46_combout ),
	.cout(\dout[13]~47 ));
defparam \dout[13]~46 .lut_mask = 16'h96BF;
defparam \dout[13]~46 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[14]~48 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4~portbdataout ),
	.datab(dout_141),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[13]~47 ),
	.combout(\dout[14]~48_combout ),
	.cout(\dout[14]~49 ));
defparam \dout[14]~48 .lut_mask = 16'h96DF;
defparam \dout[14]~48 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[15]~50 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3~portbdataout ),
	.datab(dout_151),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[14]~49 ),
	.combout(\dout[15]~50_combout ),
	.cout(\dout[15]~51 ));
defparam \dout[15]~50 .lut_mask = 16'h96BF;
defparam \dout[15]~50 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[16]~52 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2~portbdataout ),
	.datab(dout_161),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[15]~51 ),
	.combout(\dout[16]~52_combout ),
	.cout(\dout[16]~53 ));
defparam \dout[16]~52 .lut_mask = 16'h96DF;
defparam \dout[16]~52 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[17]~54 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1~portbdataout ),
	.datab(dout_171),
	.datac(gnd),
	.datad(vcc),
	.cin(\dout[16]~53 ),
	.combout(\dout[17]~54_combout ),
	.cout(\dout[17]~55 ));
defparam \dout[17]~54 .lut_mask = 16'h96BF;
defparam \dout[17]~54 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout[18]~56 (
	.dataa(\glogic:u0|register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0~portbdataout ),
	.datab(dout_181),
	.datac(gnd),
	.datad(gnd),
	.cin(\dout[17]~55 ),
	.combout(\dout[18]~56_combout ),
	.cout());
defparam \dout[18]~56 .lut_mask = 16'h9696;
defparam \dout[18]~56 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dout_valid~0 (
	.dataa(reset_n),
	.datab(dout_valid2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\dout_valid~0_combout ),
	.cout());
defparam \dout_valid~0 .lut_mask = 16'hEEEE;
defparam \dout_valid~0 .sum_lutc_input = "datac";

endmodule

module cic_auk_dspip_delay_2 (
	ram_block5a18,
	dout_0,
	ram_block5a17,
	dout_1,
	ram_block5a16,
	dout_2,
	ram_block5a15,
	dout_3,
	ram_block5a14,
	dout_4,
	ram_block5a13,
	dout_5,
	ram_block5a12,
	dout_6,
	ram_block5a11,
	dout_7,
	ram_block5a10,
	dout_8,
	ram_block5a9,
	dout_9,
	ram_block5a8,
	dout_10,
	ram_block5a7,
	dout_11,
	ram_block5a6,
	dout_12,
	ram_block5a5,
	dout_13,
	ram_block5a4,
	dout_14,
	ram_block5a3,
	dout_15,
	ram_block5a2,
	dout_16,
	ram_block5a1,
	dout_17,
	ram_block5a0,
	dout_18,
	stall_reg,
	dout_valid,
	ena_and_valid,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	ram_block5a18;
input 	dout_0;
output 	ram_block5a17;
input 	dout_1;
output 	ram_block5a16;
input 	dout_2;
output 	ram_block5a15;
input 	dout_3;
output 	ram_block5a14;
input 	dout_4;
output 	ram_block5a13;
input 	dout_5;
output 	ram_block5a12;
input 	dout_6;
output 	ram_block5a11;
input 	dout_7;
output 	ram_block5a10;
input 	dout_8;
output 	ram_block5a9;
input 	dout_9;
output 	ram_block5a8;
input 	dout_10;
output 	ram_block5a7;
input 	dout_11;
output 	ram_block5a6;
input 	dout_12;
output 	ram_block5a5;
input 	dout_13;
output 	ram_block5a4;
input 	dout_14;
output 	ram_block5a3;
input 	dout_15;
output 	ram_block5a2;
input 	dout_16;
output 	ram_block5a1;
input 	dout_17;
output 	ram_block5a0;
input 	dout_18;
input 	stall_reg;
input 	dout_valid;
input 	ena_and_valid;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0~combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[0]~q ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0~COUT ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1~combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[1]~q ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1~COUT ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~q ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~COUT ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~0_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~0_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~1 ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~2_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~3 ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~4_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~2_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~5 ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[3]~6_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual~combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0_combout ;
wire \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ;

wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1_PORTBDATAOUT_bus ;
wire [143:0] \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0_PORTBDATAOUT_bus ;

assign ram_block5a18 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18_PORTBDATAOUT_bus [0];

assign ram_block5a17 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17_PORTBDATAOUT_bus [0];

assign ram_block5a16 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16_PORTBDATAOUT_bus [0];

assign ram_block5a15 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15_PORTBDATAOUT_bus [0];

assign ram_block5a14 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14_PORTBDATAOUT_bus [0];

assign ram_block5a13 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13_PORTBDATAOUT_bus [0];

assign ram_block5a12 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12_PORTBDATAOUT_bus [0];

assign ram_block5a11 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11_PORTBDATAOUT_bus [0];

assign ram_block5a10 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10_PORTBDATAOUT_bus [0];

assign ram_block5a9 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9_PORTBDATAOUT_bus [0];

assign ram_block5a8 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8_PORTBDATAOUT_bus [0];

assign ram_block5a7 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7_PORTBDATAOUT_bus [0];

assign ram_block5a6 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6_PORTBDATAOUT_bus [0];

assign ram_block5a5 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5_PORTBDATAOUT_bus [0];

assign ram_block5a4 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4_PORTBDATAOUT_bus [0];

assign ram_block5a3 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3_PORTBDATAOUT_bus [0];

assign ram_block5a2 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2_PORTBDATAOUT_bus [0];

assign ram_block5a1 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1_PORTBDATAOUT_bus [0];

assign ram_block5a0 = \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0_PORTBDATAOUT_bus [0];

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_0}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[2].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_first_bit_number = 18;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_first_bit_number = 18;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a18 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_1}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[2].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_first_bit_number = 17;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_first_bit_number = 17;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a17 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_2}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[2].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_first_bit_number = 16;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_first_bit_number = 16;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a16 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_3}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[2].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_first_bit_number = 15;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_first_bit_number = 15;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a15 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_4}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[2].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_first_bit_number = 14;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_first_bit_number = 14;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a14 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_5}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[2].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_first_bit_number = 13;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_first_bit_number = 13;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a13 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_6}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[2].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_first_bit_number = 12;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_first_bit_number = 12;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a12 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_7}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[2].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_first_bit_number = 11;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_first_bit_number = 11;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a11 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_8}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[2].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_first_bit_number = 10;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_first_bit_number = 10;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a10 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_9}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[2].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_first_bit_number = 9;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_first_bit_number = 9;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a9 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_10}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[2].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_first_bit_number = 8;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_first_bit_number = 8;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a8 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_11}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[2].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_first_bit_number = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_first_bit_number = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a7 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_12}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[2].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_first_bit_number = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_first_bit_number = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a6 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_13}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[2].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_first_bit_number = 5;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_first_bit_number = 5;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a5 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_14}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[2].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_first_bit_number = 4;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_first_bit_number = 4;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a4 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_15}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[2].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_first_bit_number = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_first_bit_number = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a3 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_16}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[2].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_first_bit_number = 2;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_first_bit_number = 2;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a2 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_17}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[2].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_first_bit_number = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_first_bit_number = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a1 .ram_block_type = "auto";

fiftyfivenm_ram_block \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(ena_and_valid),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dout_18}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0_PORTBDATAOUT_bus ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .clk0_core_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .clk0_input_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .clk0_output_clock_enable = "ena0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .data_interleave_offset_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .data_interleave_width_in_bits = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|alt_cic_dec_miso:dec_mul|auk_dspip_differentiator:stage_diff[2].auk_dsp_diff|auk_dspip_delay:\\glogic:u0|altshift_taps:\\register_fifo:fifo_data[0][18]_rtl_0|shift_taps_qgm:auto_generated|altsyncram_6da1:altsyncram2|ALTSYNCRAM";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .mixed_port_feed_through_mode = "old";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .operation_mode = "dual_port";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_data_out_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_data_out_clock = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_first_bit_number = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_address_clear = "none";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_address_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_address_width = 3;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_data_out_clear = "clear0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_data_out_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_data_width = 1;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_first_address = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_first_bit_number = 0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_last_address = 6;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_logical_ram_depth = 7;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_logical_ram_width = 19;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .port_b_read_enable_clock = "clock0";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|altsyncram2|ram_block5a0 .ram_block_type = "auto";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0~combout ),
	.cout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0~COUT ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0 .lut_mask = 16'h55AA;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0 (
	.dataa(stall_reg),
	.datab(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~0_combout ),
	.datac(gnd),
	.datad(dout_valid),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0 .lut_mask = 16'hFF77;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0_combout ),
	.q(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[0] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita0~COUT ),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1~combout ),
	.cout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1~COUT ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1 .lut_mask = 16'h5A5F;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0_combout ),
	.q(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[1] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita1~COUT ),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~combout ),
	.cout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~COUT ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2 .lut_mask = 16'h5AAF;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~0_combout ),
	.q(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_reg_bit[2] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~COUT ),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~0_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~0 .lut_mask = 16'hF0F0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~0 .sum_lutc_input = "cin";

dffeas \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4 (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr3|counter_comb_bita2~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena_and_valid),
	.q(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4 .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|dffe4 .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~0 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~0_combout ),
	.cout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~1 ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~0 .lut_mask = 16'h55AA;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~2 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~1 ),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~2_combout ),
	.cout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~3 ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~2 .lut_mask = 16'h5A5F;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1 .lut_mask = 16'hAAFF;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena_and_valid),
	.q(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~4 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[1]~3 ),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~4_combout ),
	.cout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~5 ));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~4 .lut_mask = 16'h5AAF;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~2 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~2_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~2 .lut_mask = 16'hAAFF;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~2 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena_and_valid),
	.q(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[3]~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[2]~5 ),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[3]~6_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[3]~6 .lut_mask = 16'hF0F0;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[3]~6 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[3]~6_combout ),
	.datab(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datac(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datad(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual .lut_mask = 16'hFEFF;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0 (
	.dataa(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|add_sub6_result_int[0]~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0 .lut_mask = 16'hAAFF;
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0 .sum_lutc_input = "datac";

dffeas \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|trigger_mux_w[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena_and_valid),
	.q(\register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18]_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .power_up = "low";

endmodule

module cic_auk_dspip_downsample (
	sample_state_0,
	count_6,
	count_1,
	count_2,
	count_3,
	count_4,
	count_0,
	count_5,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	sample_state_0;
output 	count_6;
output 	count_1;
output 	count_2;
output 	count_3;
output 	count_4;
output 	count_0;
output 	count_5;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_counter_module_1 counter_fs_inst(
	.sample_state_0(sample_state_0),
	.count_6(count_6),
	.count_1(count_1),
	.count_2(count_2),
	.count_3(count_3),
	.count_4(count_4),
	.count_0(count_0),
	.count_5(count_5),
	.stall_reg(stall_reg),
	.clk(clk),
	.reset_n(reset_n));

endmodule

module cic_counter_module_1 (
	sample_state_0,
	count_6,
	count_1,
	count_2,
	count_3,
	count_4,
	count_0,
	count_5,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	sample_state_0;
output 	count_6;
output 	count_1;
output 	count_2;
output 	count_3;
output 	count_4;
output 	count_0;
output 	count_5;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \count[0]~8 ;
wire \count[1]~10 ;
wire \count[2]~12 ;
wire \count[3]~14 ;
wire \count[4]~16 ;
wire \count[5]~18 ;
wire \count[6]~19_combout ;
wire \count[1]~21_combout ;
wire \count[1]~22_combout ;
wire \count[1]~23_combout ;
wire \count[1]~24_combout ;
wire \count[1]~9_combout ;
wire \count[2]~11_combout ;
wire \count[3]~13_combout ;
wire \count[4]~15_combout ;
wire \count[0]~7_combout ;
wire \count[5]~17_combout ;


dffeas \count[6] (
	.clk(clk),
	.d(\count[6]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\count[1]~23_combout ),
	.sload(gnd),
	.ena(\count[1]~24_combout ),
	.q(count_6),
	.prn(vcc));
defparam \count[6] .is_wysiwyg = "true";
defparam \count[6] .power_up = "low";

dffeas \count[1] (
	.clk(clk),
	.d(\count[1]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\count[1]~23_combout ),
	.sload(gnd),
	.ena(\count[1]~24_combout ),
	.q(count_1),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

dffeas \count[2] (
	.clk(clk),
	.d(\count[2]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\count[1]~23_combout ),
	.sload(gnd),
	.ena(\count[1]~24_combout ),
	.q(count_2),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

dffeas \count[3] (
	.clk(clk),
	.d(\count[3]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\count[1]~23_combout ),
	.sload(gnd),
	.ena(\count[1]~24_combout ),
	.q(count_3),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

dffeas \count[4] (
	.clk(clk),
	.d(\count[4]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\count[1]~23_combout ),
	.sload(gnd),
	.ena(\count[1]~24_combout ),
	.q(count_4),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

dffeas \count[0] (
	.clk(clk),
	.d(\count[0]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\count[1]~23_combout ),
	.sload(gnd),
	.ena(\count[1]~24_combout ),
	.q(count_0),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

dffeas \count[5] (
	.clk(clk),
	.d(\count[5]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\count[1]~23_combout ),
	.sload(gnd),
	.ena(\count[1]~24_combout ),
	.q(count_5),
	.prn(vcc));
defparam \count[5] .is_wysiwyg = "true";
defparam \count[5] .power_up = "low";

fiftyfivenm_lcell_comb \count[0]~7 (
	.dataa(count_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\count[0]~7_combout ),
	.cout(\count[0]~8 ));
defparam \count[0]~7 .lut_mask = 16'h55AA;
defparam \count[0]~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \count[1]~9 (
	.dataa(count_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[0]~8 ),
	.combout(\count[1]~9_combout ),
	.cout(\count[1]~10 ));
defparam \count[1]~9 .lut_mask = 16'h5A5F;
defparam \count[1]~9 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \count[2]~11 (
	.dataa(count_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[1]~10 ),
	.combout(\count[2]~11_combout ),
	.cout(\count[2]~12 ));
defparam \count[2]~11 .lut_mask = 16'h5AAF;
defparam \count[2]~11 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \count[3]~13 (
	.dataa(count_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[2]~12 ),
	.combout(\count[3]~13_combout ),
	.cout(\count[3]~14 ));
defparam \count[3]~13 .lut_mask = 16'h5A5F;
defparam \count[3]~13 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \count[4]~15 (
	.dataa(count_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[3]~14 ),
	.combout(\count[4]~15_combout ),
	.cout(\count[4]~16 ));
defparam \count[4]~15 .lut_mask = 16'h5AAF;
defparam \count[4]~15 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \count[5]~17 (
	.dataa(count_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\count[4]~16 ),
	.combout(\count[5]~17_combout ),
	.cout(\count[5]~18 ));
defparam \count[5]~17 .lut_mask = 16'h5A5F;
defparam \count[5]~17 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \count[6]~19 (
	.dataa(count_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\count[5]~18 ),
	.combout(\count[6]~19_combout ),
	.cout());
defparam \count[6]~19 .lut_mask = 16'h5A5A;
defparam \count[6]~19 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \count[1]~21 (
	.dataa(count_0),
	.datab(count_1),
	.datac(count_2),
	.datad(count_3),
	.cin(gnd),
	.combout(\count[1]~21_combout ),
	.cout());
defparam \count[1]~21 .lut_mask = 16'h7FFF;
defparam \count[1]~21 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \count[1]~22 (
	.dataa(count_6),
	.datab(gnd),
	.datac(count_5),
	.datad(count_4),
	.cin(gnd),
	.combout(\count[1]~22_combout ),
	.cout());
defparam \count[1]~22 .lut_mask = 16'hAFFF;
defparam \count[1]~22 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \count[1]~23 (
	.dataa(reset_n),
	.datab(\count[1]~21_combout ),
	.datac(\count[1]~22_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\count[1]~23_combout ),
	.cout());
defparam \count[1]~23 .lut_mask = 16'h7F7F;
defparam \count[1]~23 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \count[1]~24 (
	.dataa(reset_n),
	.datab(stall_reg),
	.datac(gnd),
	.datad(sample_state_0),
	.cin(gnd),
	.combout(\count[1]~24_combout ),
	.cout());
defparam \count[1]~24 .lut_mask = 16'hFF77;
defparam \count[1]~24 .sum_lutc_input = "datac";

endmodule

module cic_auk_dspip_integrator (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	q_b_0,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	q_b_0;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_3 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.q_b_0(q_b_0),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_3 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	q_b_0,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	q_b_0;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(q_b_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(q_b_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(q_b_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(q_b_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(q_b_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_0),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_0),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_1 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_4 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data001(register_fifofifo_data001),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data051(register_fifofifo_data051),
	.register_fifofifo_data061(register_fifofifo_data061),
	.register_fifofifo_data071(register_fifofifo_data071),
	.register_fifofifo_data081(register_fifofifo_data081),
	.register_fifofifo_data091(register_fifofifo_data091),
	.register_fifofifo_data0101(register_fifofifo_data0101),
	.register_fifofifo_data0111(register_fifofifo_data0111),
	.register_fifofifo_data0121(register_fifofifo_data0121),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.register_fifofifo_data0141(register_fifofifo_data0141),
	.register_fifofifo_data0151(register_fifofifo_data0151),
	.register_fifofifo_data0161(register_fifofifo_data0161),
	.register_fifofifo_data0171(register_fifofifo_data0171),
	.register_fifofifo_data0181(register_fifofifo_data0181),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_4 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(register_fifofifo_data001),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(register_fifofifo_data019),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(register_fifofifo_data021),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(register_fifofifo_data031),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(register_fifofifo_data041),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(register_fifofifo_data051),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(register_fifofifo_data061),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(register_fifofifo_data071),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(register_fifofifo_data081),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(register_fifofifo_data091),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(register_fifofifo_data0101),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(register_fifofifo_data0111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(register_fifofifo_data0121),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(register_fifofifo_data0131),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(register_fifofifo_data0141),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(register_fifofifo_data0151),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(register_fifofifo_data0161),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(register_fifofifo_data0171),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(register_fifofifo_data0181),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_2 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_5 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data001(register_fifofifo_data001),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data051(register_fifofifo_data051),
	.register_fifofifo_data061(register_fifofifo_data061),
	.register_fifofifo_data071(register_fifofifo_data071),
	.register_fifofifo_data081(register_fifofifo_data081),
	.register_fifofifo_data091(register_fifofifo_data091),
	.register_fifofifo_data0101(register_fifofifo_data0101),
	.register_fifofifo_data0111(register_fifofifo_data0111),
	.register_fifofifo_data0121(register_fifofifo_data0121),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.register_fifofifo_data0141(register_fifofifo_data0141),
	.register_fifofifo_data0151(register_fifofifo_data0151),
	.register_fifofifo_data0161(register_fifofifo_data0161),
	.register_fifofifo_data0171(register_fifofifo_data0171),
	.register_fifofifo_data0181(register_fifofifo_data0181),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_5 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(register_fifofifo_data001),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(register_fifofifo_data019),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(register_fifofifo_data021),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(register_fifofifo_data031),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(register_fifofifo_data041),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(register_fifofifo_data051),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(register_fifofifo_data061),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(register_fifofifo_data071),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(register_fifofifo_data081),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(register_fifofifo_data091),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(register_fifofifo_data0101),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(register_fifofifo_data0111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(register_fifofifo_data0121),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(register_fifofifo_data0131),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(register_fifofifo_data0141),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(register_fifofifo_data0151),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(register_fifofifo_data0161),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(register_fifofifo_data0171),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(register_fifofifo_data0181),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_3 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	q_b_1,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	q_b_1;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_6 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.q_b_1(q_b_1),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_6 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	q_b_1,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	q_b_1;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(q_b_1),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(q_b_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(q_b_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(q_b_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(q_b_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_1),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_4 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_7 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data001(register_fifofifo_data001),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data051(register_fifofifo_data051),
	.register_fifofifo_data061(register_fifofifo_data061),
	.register_fifofifo_data071(register_fifofifo_data071),
	.register_fifofifo_data081(register_fifofifo_data081),
	.register_fifofifo_data091(register_fifofifo_data091),
	.register_fifofifo_data0101(register_fifofifo_data0101),
	.register_fifofifo_data0111(register_fifofifo_data0111),
	.register_fifofifo_data0121(register_fifofifo_data0121),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.register_fifofifo_data0141(register_fifofifo_data0141),
	.register_fifofifo_data0151(register_fifofifo_data0151),
	.register_fifofifo_data0161(register_fifofifo_data0161),
	.register_fifofifo_data0171(register_fifofifo_data0171),
	.register_fifofifo_data0181(register_fifofifo_data0181),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_7 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(register_fifofifo_data001),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(register_fifofifo_data019),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(register_fifofifo_data021),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(register_fifofifo_data031),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(register_fifofifo_data041),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(register_fifofifo_data051),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(register_fifofifo_data061),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(register_fifofifo_data071),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(register_fifofifo_data081),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(register_fifofifo_data091),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(register_fifofifo_data0101),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(register_fifofifo_data0111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(register_fifofifo_data0121),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(register_fifofifo_data0131),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(register_fifofifo_data0141),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(register_fifofifo_data0151),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(register_fifofifo_data0161),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(register_fifofifo_data0171),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(register_fifofifo_data0181),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_5 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_8 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data001(register_fifofifo_data001),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data051(register_fifofifo_data051),
	.register_fifofifo_data061(register_fifofifo_data061),
	.register_fifofifo_data071(register_fifofifo_data071),
	.register_fifofifo_data081(register_fifofifo_data081),
	.register_fifofifo_data091(register_fifofifo_data091),
	.register_fifofifo_data0101(register_fifofifo_data0101),
	.register_fifofifo_data0111(register_fifofifo_data0111),
	.register_fifofifo_data0121(register_fifofifo_data0121),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.register_fifofifo_data0141(register_fifofifo_data0141),
	.register_fifofifo_data0151(register_fifofifo_data0151),
	.register_fifofifo_data0161(register_fifofifo_data0161),
	.register_fifofifo_data0171(register_fifofifo_data0171),
	.register_fifofifo_data0181(register_fifofifo_data0181),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_8 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(register_fifofifo_data001),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(register_fifofifo_data019),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(register_fifofifo_data021),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(register_fifofifo_data031),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(register_fifofifo_data041),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(register_fifofifo_data051),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(register_fifofifo_data061),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(register_fifofifo_data071),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(register_fifofifo_data081),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(register_fifofifo_data091),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(register_fifofifo_data0101),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(register_fifofifo_data0111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(register_fifofifo_data0121),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(register_fifofifo_data0131),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(register_fifofifo_data0141),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(register_fifofifo_data0151),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(register_fifofifo_data0161),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(register_fifofifo_data0171),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(register_fifofifo_data0181),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_6 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	q_b_2,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	q_b_2;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_9 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.q_b_2(q_b_2),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_9 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	q_b_2,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	q_b_2;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(q_b_2),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(q_b_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(q_b_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(q_b_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(q_b_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_2),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_7 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_10 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data001(register_fifofifo_data001),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data051(register_fifofifo_data051),
	.register_fifofifo_data061(register_fifofifo_data061),
	.register_fifofifo_data071(register_fifofifo_data071),
	.register_fifofifo_data081(register_fifofifo_data081),
	.register_fifofifo_data091(register_fifofifo_data091),
	.register_fifofifo_data0101(register_fifofifo_data0101),
	.register_fifofifo_data0111(register_fifofifo_data0111),
	.register_fifofifo_data0121(register_fifofifo_data0121),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.register_fifofifo_data0141(register_fifofifo_data0141),
	.register_fifofifo_data0151(register_fifofifo_data0151),
	.register_fifofifo_data0161(register_fifofifo_data0161),
	.register_fifofifo_data0171(register_fifofifo_data0171),
	.register_fifofifo_data0181(register_fifofifo_data0181),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_10 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(register_fifofifo_data001),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(register_fifofifo_data019),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(register_fifofifo_data021),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(register_fifofifo_data031),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(register_fifofifo_data041),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(register_fifofifo_data051),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(register_fifofifo_data061),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(register_fifofifo_data071),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(register_fifofifo_data081),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(register_fifofifo_data091),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(register_fifofifo_data0101),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(register_fifofifo_data0111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(register_fifofifo_data0121),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(register_fifofifo_data0131),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(register_fifofifo_data0141),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(register_fifofifo_data0151),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(register_fifofifo_data0161),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(register_fifofifo_data0171),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(register_fifofifo_data0181),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_8 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_11 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data001(register_fifofifo_data001),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data051(register_fifofifo_data051),
	.register_fifofifo_data061(register_fifofifo_data061),
	.register_fifofifo_data071(register_fifofifo_data071),
	.register_fifofifo_data081(register_fifofifo_data081),
	.register_fifofifo_data091(register_fifofifo_data091),
	.register_fifofifo_data0101(register_fifofifo_data0101),
	.register_fifofifo_data0111(register_fifofifo_data0111),
	.register_fifofifo_data0121(register_fifofifo_data0121),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.register_fifofifo_data0141(register_fifofifo_data0141),
	.register_fifofifo_data0151(register_fifofifo_data0151),
	.register_fifofifo_data0161(register_fifofifo_data0161),
	.register_fifofifo_data0171(register_fifofifo_data0171),
	.register_fifofifo_data0181(register_fifofifo_data0181),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_11 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(register_fifofifo_data001),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(register_fifofifo_data019),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(register_fifofifo_data021),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(register_fifofifo_data031),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(register_fifofifo_data041),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(register_fifofifo_data051),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(register_fifofifo_data061),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(register_fifofifo_data071),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(register_fifofifo_data081),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(register_fifofifo_data091),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(register_fifofifo_data0101),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(register_fifofifo_data0111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(register_fifofifo_data0121),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(register_fifofifo_data0131),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(register_fifofifo_data0141),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(register_fifofifo_data0151),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(register_fifofifo_data0161),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(register_fifofifo_data0171),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(register_fifofifo_data0181),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_9 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	q_b_3,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	q_b_3;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_12 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.q_b_3(q_b_3),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_12 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	q_b_3,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	q_b_3;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(q_b_3),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(q_b_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(q_b_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(q_b_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(q_b_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_3),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_10 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_13 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data001(register_fifofifo_data001),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data051(register_fifofifo_data051),
	.register_fifofifo_data061(register_fifofifo_data061),
	.register_fifofifo_data071(register_fifofifo_data071),
	.register_fifofifo_data081(register_fifofifo_data081),
	.register_fifofifo_data091(register_fifofifo_data091),
	.register_fifofifo_data0101(register_fifofifo_data0101),
	.register_fifofifo_data0111(register_fifofifo_data0111),
	.register_fifofifo_data0121(register_fifofifo_data0121),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.register_fifofifo_data0141(register_fifofifo_data0141),
	.register_fifofifo_data0151(register_fifofifo_data0151),
	.register_fifofifo_data0161(register_fifofifo_data0161),
	.register_fifofifo_data0171(register_fifofifo_data0171),
	.register_fifofifo_data0181(register_fifofifo_data0181),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_13 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(register_fifofifo_data001),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(register_fifofifo_data019),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(register_fifofifo_data021),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(register_fifofifo_data031),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(register_fifofifo_data041),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(register_fifofifo_data051),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(register_fifofifo_data061),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(register_fifofifo_data071),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(register_fifofifo_data081),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(register_fifofifo_data091),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(register_fifofifo_data0101),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(register_fifofifo_data0111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(register_fifofifo_data0121),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(register_fifofifo_data0131),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(register_fifofifo_data0141),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(register_fifofifo_data0151),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(register_fifofifo_data0161),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(register_fifofifo_data0171),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(register_fifofifo_data0181),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_11 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_14 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data001(register_fifofifo_data001),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data051(register_fifofifo_data051),
	.register_fifofifo_data061(register_fifofifo_data061),
	.register_fifofifo_data071(register_fifofifo_data071),
	.register_fifofifo_data081(register_fifofifo_data081),
	.register_fifofifo_data091(register_fifofifo_data091),
	.register_fifofifo_data0101(register_fifofifo_data0101),
	.register_fifofifo_data0111(register_fifofifo_data0111),
	.register_fifofifo_data0121(register_fifofifo_data0121),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.register_fifofifo_data0141(register_fifofifo_data0141),
	.register_fifofifo_data0151(register_fifofifo_data0151),
	.register_fifofifo_data0161(register_fifofifo_data0161),
	.register_fifofifo_data0171(register_fifofifo_data0171),
	.register_fifofifo_data0181(register_fifofifo_data0181),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_14 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(register_fifofifo_data001),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(register_fifofifo_data019),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(register_fifofifo_data021),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(register_fifofifo_data031),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(register_fifofifo_data041),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(register_fifofifo_data051),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(register_fifofifo_data061),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(register_fifofifo_data071),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(register_fifofifo_data081),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(register_fifofifo_data091),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(register_fifofifo_data0101),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(register_fifofifo_data0111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(register_fifofifo_data0121),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(register_fifofifo_data0131),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(register_fifofifo_data0141),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(register_fifofifo_data0151),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(register_fifofifo_data0161),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(register_fifofifo_data0171),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(register_fifofifo_data0181),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_12 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	q_b_4,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	q_b_4;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_15 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.q_b_4(q_b_4),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_15 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	q_b_4,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	q_b_4;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(q_b_4),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(q_b_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(q_b_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(q_b_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(q_b_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_4),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_13 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_16 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data001(register_fifofifo_data001),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data051(register_fifofifo_data051),
	.register_fifofifo_data061(register_fifofifo_data061),
	.register_fifofifo_data071(register_fifofifo_data071),
	.register_fifofifo_data081(register_fifofifo_data081),
	.register_fifofifo_data091(register_fifofifo_data091),
	.register_fifofifo_data0101(register_fifofifo_data0101),
	.register_fifofifo_data0111(register_fifofifo_data0111),
	.register_fifofifo_data0121(register_fifofifo_data0121),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.register_fifofifo_data0141(register_fifofifo_data0141),
	.register_fifofifo_data0151(register_fifofifo_data0151),
	.register_fifofifo_data0161(register_fifofifo_data0161),
	.register_fifofifo_data0171(register_fifofifo_data0171),
	.register_fifofifo_data0181(register_fifofifo_data0181),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_16 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(register_fifofifo_data001),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(register_fifofifo_data019),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(register_fifofifo_data021),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(register_fifofifo_data031),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(register_fifofifo_data041),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(register_fifofifo_data051),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(register_fifofifo_data061),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(register_fifofifo_data071),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(register_fifofifo_data081),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(register_fifofifo_data091),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(register_fifofifo_data0101),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(register_fifofifo_data0111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(register_fifofifo_data0121),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(register_fifofifo_data0131),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(register_fifofifo_data0141),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(register_fifofifo_data0151),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(register_fifofifo_data0161),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(register_fifofifo_data0171),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(register_fifofifo_data0181),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_14 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_17 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data001(register_fifofifo_data001),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data051(register_fifofifo_data051),
	.register_fifofifo_data061(register_fifofifo_data061),
	.register_fifofifo_data071(register_fifofifo_data071),
	.register_fifofifo_data081(register_fifofifo_data081),
	.register_fifofifo_data091(register_fifofifo_data091),
	.register_fifofifo_data0101(register_fifofifo_data0101),
	.register_fifofifo_data0111(register_fifofifo_data0111),
	.register_fifofifo_data0121(register_fifofifo_data0121),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.register_fifofifo_data0141(register_fifofifo_data0141),
	.register_fifofifo_data0151(register_fifofifo_data0151),
	.register_fifofifo_data0161(register_fifofifo_data0161),
	.register_fifofifo_data0171(register_fifofifo_data0171),
	.register_fifofifo_data0181(register_fifofifo_data0181),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_17 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(register_fifofifo_data001),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(register_fifofifo_data019),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(register_fifofifo_data021),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(register_fifofifo_data031),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(register_fifofifo_data041),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(register_fifofifo_data051),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(register_fifofifo_data061),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(register_fifofifo_data071),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(register_fifofifo_data081),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(register_fifofifo_data091),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(register_fifofifo_data0101),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(register_fifofifo_data0111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(register_fifofifo_data0121),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(register_fifofifo_data0131),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(register_fifofifo_data0141),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(register_fifofifo_data0151),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(register_fifofifo_data0161),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(register_fifofifo_data0171),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(register_fifofifo_data0181),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_15 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	q_b_5,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	q_b_5;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_18 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.q_b_5(q_b_5),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_18 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	q_b_5,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	q_b_5;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(q_b_5),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(q_b_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(q_b_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(q_b_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(q_b_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_5),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_16 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_19 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data001(register_fifofifo_data001),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data051(register_fifofifo_data051),
	.register_fifofifo_data061(register_fifofifo_data061),
	.register_fifofifo_data071(register_fifofifo_data071),
	.register_fifofifo_data081(register_fifofifo_data081),
	.register_fifofifo_data091(register_fifofifo_data091),
	.register_fifofifo_data0101(register_fifofifo_data0101),
	.register_fifofifo_data0111(register_fifofifo_data0111),
	.register_fifofifo_data0121(register_fifofifo_data0121),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.register_fifofifo_data0141(register_fifofifo_data0141),
	.register_fifofifo_data0151(register_fifofifo_data0151),
	.register_fifofifo_data0161(register_fifofifo_data0161),
	.register_fifofifo_data0171(register_fifofifo_data0171),
	.register_fifofifo_data0181(register_fifofifo_data0181),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_19 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(register_fifofifo_data001),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(register_fifofifo_data019),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(register_fifofifo_data021),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(register_fifofifo_data031),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(register_fifofifo_data041),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(register_fifofifo_data051),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(register_fifofifo_data061),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(register_fifofifo_data071),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(register_fifofifo_data081),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(register_fifofifo_data091),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(register_fifofifo_data0101),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(register_fifofifo_data0111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(register_fifofifo_data0121),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(register_fifofifo_data0131),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(register_fifofifo_data0141),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(register_fifofifo_data0151),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(register_fifofifo_data0161),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(register_fifofifo_data0171),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(register_fifofifo_data0181),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_17 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_20 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data001(register_fifofifo_data001),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data051(register_fifofifo_data051),
	.register_fifofifo_data061(register_fifofifo_data061),
	.register_fifofifo_data071(register_fifofifo_data071),
	.register_fifofifo_data081(register_fifofifo_data081),
	.register_fifofifo_data091(register_fifofifo_data091),
	.register_fifofifo_data0101(register_fifofifo_data0101),
	.register_fifofifo_data0111(register_fifofifo_data0111),
	.register_fifofifo_data0121(register_fifofifo_data0121),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.register_fifofifo_data0141(register_fifofifo_data0141),
	.register_fifofifo_data0151(register_fifofifo_data0151),
	.register_fifofifo_data0161(register_fifofifo_data0161),
	.register_fifofifo_data0171(register_fifofifo_data0171),
	.register_fifofifo_data0181(register_fifofifo_data0181),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_20 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(register_fifofifo_data001),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(register_fifofifo_data019),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(register_fifofifo_data021),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(register_fifofifo_data031),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(register_fifofifo_data041),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(register_fifofifo_data051),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(register_fifofifo_data061),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(register_fifofifo_data071),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(register_fifofifo_data081),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(register_fifofifo_data091),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(register_fifofifo_data0101),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(register_fifofifo_data0111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(register_fifofifo_data0121),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(register_fifofifo_data0131),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(register_fifofifo_data0141),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(register_fifofifo_data0151),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(register_fifofifo_data0161),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(register_fifofifo_data0171),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(register_fifofifo_data0181),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_18 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	q_b_6,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	q_b_6;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_21 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.q_b_6(q_b_6),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_21 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	q_b_6,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	q_b_6;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(q_b_6),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(q_b_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(q_b_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(q_b_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(q_b_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_6),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_19 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_22 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data001(register_fifofifo_data001),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data051(register_fifofifo_data051),
	.register_fifofifo_data061(register_fifofifo_data061),
	.register_fifofifo_data071(register_fifofifo_data071),
	.register_fifofifo_data081(register_fifofifo_data081),
	.register_fifofifo_data091(register_fifofifo_data091),
	.register_fifofifo_data0101(register_fifofifo_data0101),
	.register_fifofifo_data0111(register_fifofifo_data0111),
	.register_fifofifo_data0121(register_fifofifo_data0121),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.register_fifofifo_data0141(register_fifofifo_data0141),
	.register_fifofifo_data0151(register_fifofifo_data0151),
	.register_fifofifo_data0161(register_fifofifo_data0161),
	.register_fifofifo_data0171(register_fifofifo_data0171),
	.register_fifofifo_data0181(register_fifofifo_data0181),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_22 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(register_fifofifo_data001),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(register_fifofifo_data019),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(register_fifofifo_data021),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(register_fifofifo_data031),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(register_fifofifo_data041),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(register_fifofifo_data051),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(register_fifofifo_data061),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(register_fifofifo_data071),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(register_fifofifo_data081),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(register_fifofifo_data091),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(register_fifofifo_data0101),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(register_fifofifo_data0111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(register_fifofifo_data0121),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(register_fifofifo_data0131),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(register_fifofifo_data0141),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(register_fifofifo_data0151),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(register_fifofifo_data0161),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(register_fifofifo_data0171),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(register_fifofifo_data0181),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_20 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_23 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data001(register_fifofifo_data001),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data051(register_fifofifo_data051),
	.register_fifofifo_data061(register_fifofifo_data061),
	.register_fifofifo_data071(register_fifofifo_data071),
	.register_fifofifo_data081(register_fifofifo_data081),
	.register_fifofifo_data091(register_fifofifo_data091),
	.register_fifofifo_data0101(register_fifofifo_data0101),
	.register_fifofifo_data0111(register_fifofifo_data0111),
	.register_fifofifo_data0121(register_fifofifo_data0121),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.register_fifofifo_data0141(register_fifofifo_data0141),
	.register_fifofifo_data0151(register_fifofifo_data0151),
	.register_fifofifo_data0161(register_fifofifo_data0161),
	.register_fifofifo_data0171(register_fifofifo_data0171),
	.register_fifofifo_data0181(register_fifofifo_data0181),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_23 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(register_fifofifo_data001),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(register_fifofifo_data019),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(register_fifofifo_data021),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(register_fifofifo_data031),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(register_fifofifo_data041),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(register_fifofifo_data051),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(register_fifofifo_data061),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(register_fifofifo_data071),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(register_fifofifo_data081),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(register_fifofifo_data091),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(register_fifofifo_data0101),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(register_fifofifo_data0111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(register_fifofifo_data0121),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(register_fifofifo_data0131),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(register_fifofifo_data0141),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(register_fifofifo_data0151),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(register_fifofifo_data0161),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(register_fifofifo_data0171),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(register_fifofifo_data0181),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_21 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	q_b_7,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	q_b_7;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_24 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.q_b_7(q_b_7),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_24 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	q_b_7,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	q_b_7;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(q_b_7),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(q_b_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(q_b_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(q_b_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(q_b_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_7),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_22 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_25 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data001(register_fifofifo_data001),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data051(register_fifofifo_data051),
	.register_fifofifo_data061(register_fifofifo_data061),
	.register_fifofifo_data071(register_fifofifo_data071),
	.register_fifofifo_data081(register_fifofifo_data081),
	.register_fifofifo_data091(register_fifofifo_data091),
	.register_fifofifo_data0101(register_fifofifo_data0101),
	.register_fifofifo_data0111(register_fifofifo_data0111),
	.register_fifofifo_data0121(register_fifofifo_data0121),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.register_fifofifo_data0141(register_fifofifo_data0141),
	.register_fifofifo_data0151(register_fifofifo_data0151),
	.register_fifofifo_data0161(register_fifofifo_data0161),
	.register_fifofifo_data0171(register_fifofifo_data0171),
	.register_fifofifo_data0181(register_fifofifo_data0181),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_25 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(register_fifofifo_data001),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(register_fifofifo_data019),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(register_fifofifo_data021),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(register_fifofifo_data031),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(register_fifofifo_data041),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(register_fifofifo_data051),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(register_fifofifo_data061),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(register_fifofifo_data071),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(register_fifofifo_data081),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(register_fifofifo_data091),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(register_fifofifo_data0101),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(register_fifofifo_data0111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(register_fifofifo_data0121),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(register_fifofifo_data0131),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(register_fifofifo_data0141),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(register_fifofifo_data0151),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(register_fifofifo_data0161),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(register_fifofifo_data0171),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(register_fifofifo_data0181),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_23 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_26 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data001(register_fifofifo_data001),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data051(register_fifofifo_data051),
	.register_fifofifo_data061(register_fifofifo_data061),
	.register_fifofifo_data071(register_fifofifo_data071),
	.register_fifofifo_data081(register_fifofifo_data081),
	.register_fifofifo_data091(register_fifofifo_data091),
	.register_fifofifo_data0101(register_fifofifo_data0101),
	.register_fifofifo_data0111(register_fifofifo_data0111),
	.register_fifofifo_data0121(register_fifofifo_data0121),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.register_fifofifo_data0141(register_fifofifo_data0141),
	.register_fifofifo_data0151(register_fifofifo_data0151),
	.register_fifofifo_data0161(register_fifofifo_data0161),
	.register_fifofifo_data0171(register_fifofifo_data0171),
	.register_fifofifo_data0181(register_fifofifo_data0181),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_26 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(register_fifofifo_data001),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(register_fifofifo_data019),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(register_fifofifo_data021),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(register_fifofifo_data031),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(register_fifofifo_data041),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(register_fifofifo_data051),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(register_fifofifo_data061),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(register_fifofifo_data071),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(register_fifofifo_data081),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(register_fifofifo_data091),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(register_fifofifo_data0101),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(register_fifofifo_data0111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(register_fifofifo_data0121),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(register_fifofifo_data0131),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(register_fifofifo_data0141),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(register_fifofifo_data0151),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(register_fifofifo_data0161),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(register_fifofifo_data0171),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(register_fifofifo_data0181),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_24 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	q_b_8,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	q_b_8;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_27 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.q_b_8(q_b_8),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_27 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	q_b_8,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	q_b_8;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(q_b_8),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(q_b_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(q_b_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(q_b_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(q_b_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(q_b_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(q_b_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(q_b_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(q_b_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(q_b_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(q_b_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(q_b_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(q_b_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(q_b_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(q_b_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(q_b_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(q_b_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(q_b_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(q_b_8),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_25 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_28 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data001(register_fifofifo_data001),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data051(register_fifofifo_data051),
	.register_fifofifo_data061(register_fifofifo_data061),
	.register_fifofifo_data071(register_fifofifo_data071),
	.register_fifofifo_data081(register_fifofifo_data081),
	.register_fifofifo_data091(register_fifofifo_data091),
	.register_fifofifo_data0101(register_fifofifo_data0101),
	.register_fifofifo_data0111(register_fifofifo_data0111),
	.register_fifofifo_data0121(register_fifofifo_data0121),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.register_fifofifo_data0141(register_fifofifo_data0141),
	.register_fifofifo_data0151(register_fifofifo_data0151),
	.register_fifofifo_data0161(register_fifofifo_data0161),
	.register_fifofifo_data0171(register_fifofifo_data0171),
	.register_fifofifo_data0181(register_fifofifo_data0181),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_28 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(register_fifofifo_data001),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(register_fifofifo_data019),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(register_fifofifo_data021),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(register_fifofifo_data031),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(register_fifofifo_data041),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(register_fifofifo_data051),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(register_fifofifo_data061),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(register_fifofifo_data071),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(register_fifofifo_data081),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(register_fifofifo_data091),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(register_fifofifo_data0101),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(register_fifofifo_data0111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(register_fifofifo_data0121),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(register_fifofifo_data0131),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(register_fifofifo_data0141),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(register_fifofifo_data0151),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(register_fifofifo_data0161),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(register_fifofifo_data0171),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(register_fifofifo_data0181),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_auk_dspip_integrator_26 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	stall_reg,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	stall_reg;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_auk_dspip_delay_29 \glogic:integrator_pipeline_0_generate:u1 (
	.register_fifofifo_data00(register_fifofifo_data00),
	.register_fifofifo_data01(register_fifofifo_data01),
	.register_fifofifo_data02(register_fifofifo_data02),
	.register_fifofifo_data03(register_fifofifo_data03),
	.register_fifofifo_data04(register_fifofifo_data04),
	.register_fifofifo_data05(register_fifofifo_data05),
	.register_fifofifo_data06(register_fifofifo_data06),
	.register_fifofifo_data07(register_fifofifo_data07),
	.register_fifofifo_data08(register_fifofifo_data08),
	.register_fifofifo_data09(register_fifofifo_data09),
	.register_fifofifo_data010(register_fifofifo_data010),
	.register_fifofifo_data011(register_fifofifo_data011),
	.register_fifofifo_data012(register_fifofifo_data012),
	.register_fifofifo_data013(register_fifofifo_data013),
	.register_fifofifo_data014(register_fifofifo_data014),
	.register_fifofifo_data015(register_fifofifo_data015),
	.register_fifofifo_data016(register_fifofifo_data016),
	.register_fifofifo_data017(register_fifofifo_data017),
	.register_fifofifo_data018(register_fifofifo_data018),
	.register_fifofifo_data001(register_fifofifo_data001),
	.register_fifofifo_data019(register_fifofifo_data019),
	.register_fifofifo_data021(register_fifofifo_data021),
	.register_fifofifo_data031(register_fifofifo_data031),
	.register_fifofifo_data041(register_fifofifo_data041),
	.register_fifofifo_data051(register_fifofifo_data051),
	.register_fifofifo_data061(register_fifofifo_data061),
	.register_fifofifo_data071(register_fifofifo_data071),
	.register_fifofifo_data081(register_fifofifo_data081),
	.register_fifofifo_data091(register_fifofifo_data091),
	.register_fifofifo_data0101(register_fifofifo_data0101),
	.register_fifofifo_data0111(register_fifofifo_data0111),
	.register_fifofifo_data0121(register_fifofifo_data0121),
	.register_fifofifo_data0131(register_fifofifo_data0131),
	.register_fifofifo_data0141(register_fifofifo_data0141),
	.register_fifofifo_data0151(register_fifofifo_data0151),
	.register_fifofifo_data0161(register_fifofifo_data0161),
	.register_fifofifo_data0171(register_fifofifo_data0171),
	.register_fifofifo_data0181(register_fifofifo_data0181),
	.enable(stall_reg),
	.clk(clk),
	.reset(reset_n));

endmodule

module cic_auk_dspip_delay_29 (
	register_fifofifo_data00,
	register_fifofifo_data01,
	register_fifofifo_data02,
	register_fifofifo_data03,
	register_fifofifo_data04,
	register_fifofifo_data05,
	register_fifofifo_data06,
	register_fifofifo_data07,
	register_fifofifo_data08,
	register_fifofifo_data09,
	register_fifofifo_data010,
	register_fifofifo_data011,
	register_fifofifo_data012,
	register_fifofifo_data013,
	register_fifofifo_data014,
	register_fifofifo_data015,
	register_fifofifo_data016,
	register_fifofifo_data017,
	register_fifofifo_data018,
	register_fifofifo_data001,
	register_fifofifo_data019,
	register_fifofifo_data021,
	register_fifofifo_data031,
	register_fifofifo_data041,
	register_fifofifo_data051,
	register_fifofifo_data061,
	register_fifofifo_data071,
	register_fifofifo_data081,
	register_fifofifo_data091,
	register_fifofifo_data0101,
	register_fifofifo_data0111,
	register_fifofifo_data0121,
	register_fifofifo_data0131,
	register_fifofifo_data0141,
	register_fifofifo_data0151,
	register_fifofifo_data0161,
	register_fifofifo_data0171,
	register_fifofifo_data0181,
	enable,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	register_fifofifo_data00;
output 	register_fifofifo_data01;
output 	register_fifofifo_data02;
output 	register_fifofifo_data03;
output 	register_fifofifo_data04;
output 	register_fifofifo_data05;
output 	register_fifofifo_data06;
output 	register_fifofifo_data07;
output 	register_fifofifo_data08;
output 	register_fifofifo_data09;
output 	register_fifofifo_data010;
output 	register_fifofifo_data011;
output 	register_fifofifo_data012;
output 	register_fifofifo_data013;
output 	register_fifofifo_data014;
output 	register_fifofifo_data015;
output 	register_fifofifo_data016;
output 	register_fifofifo_data017;
output 	register_fifofifo_data018;
input 	register_fifofifo_data001;
input 	register_fifofifo_data019;
input 	register_fifofifo_data021;
input 	register_fifofifo_data031;
input 	register_fifofifo_data041;
input 	register_fifofifo_data051;
input 	register_fifofifo_data061;
input 	register_fifofifo_data071;
input 	register_fifofifo_data081;
input 	register_fifofifo_data091;
input 	register_fifofifo_data0101;
input 	register_fifofifo_data0111;
input 	register_fifofifo_data0121;
input 	register_fifofifo_data0131;
input 	register_fifofifo_data0141;
input 	register_fifofifo_data0151;
input 	register_fifofifo_data0161;
input 	register_fifofifo_data0171;
input 	register_fifofifo_data0181;
input 	enable;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \register_fifo:fifo_data[0][0]~1_combout ;
wire \register_fifo:fifo_data[0][0]~2 ;
wire \register_fifo:fifo_data[0][1]~1_combout ;
wire \register_fifo:fifo_data[0][1]~2 ;
wire \register_fifo:fifo_data[0][2]~1_combout ;
wire \register_fifo:fifo_data[0][2]~2 ;
wire \register_fifo:fifo_data[0][3]~1_combout ;
wire \register_fifo:fifo_data[0][3]~2 ;
wire \register_fifo:fifo_data[0][4]~1_combout ;
wire \register_fifo:fifo_data[0][4]~2 ;
wire \register_fifo:fifo_data[0][5]~1_combout ;
wire \register_fifo:fifo_data[0][5]~2 ;
wire \register_fifo:fifo_data[0][6]~1_combout ;
wire \register_fifo:fifo_data[0][6]~2 ;
wire \register_fifo:fifo_data[0][7]~1_combout ;
wire \register_fifo:fifo_data[0][7]~2 ;
wire \register_fifo:fifo_data[0][8]~1_combout ;
wire \register_fifo:fifo_data[0][8]~2 ;
wire \register_fifo:fifo_data[0][9]~1_combout ;
wire \register_fifo:fifo_data[0][9]~2 ;
wire \register_fifo:fifo_data[0][10]~1_combout ;
wire \register_fifo:fifo_data[0][10]~2 ;
wire \register_fifo:fifo_data[0][11]~1_combout ;
wire \register_fifo:fifo_data[0][11]~2 ;
wire \register_fifo:fifo_data[0][12]~1_combout ;
wire \register_fifo:fifo_data[0][12]~2 ;
wire \register_fifo:fifo_data[0][13]~1_combout ;
wire \register_fifo:fifo_data[0][13]~2 ;
wire \register_fifo:fifo_data[0][14]~1_combout ;
wire \register_fifo:fifo_data[0][14]~2 ;
wire \register_fifo:fifo_data[0][15]~1_combout ;
wire \register_fifo:fifo_data[0][15]~2 ;
wire \register_fifo:fifo_data[0][16]~1_combout ;
wire \register_fifo:fifo_data[0][16]~2 ;
wire \register_fifo:fifo_data[0][17]~1_combout ;
wire \register_fifo:fifo_data[0][17]~2 ;
wire \register_fifo:fifo_data[0][18]~1_combout ;


dffeas \register_fifo:fifo_data[0][0] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data00),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][0] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][0] .power_up = "low";

dffeas \register_fifo:fifo_data[0][1] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data01),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][1] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][1] .power_up = "low";

dffeas \register_fifo:fifo_data[0][2] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data02),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][2] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][2] .power_up = "low";

dffeas \register_fifo:fifo_data[0][3] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data03),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][3] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][3] .power_up = "low";

dffeas \register_fifo:fifo_data[0][4] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][4]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data04),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][4] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][4] .power_up = "low";

dffeas \register_fifo:fifo_data[0][5] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][5]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data05),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][5] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][5] .power_up = "low";

dffeas \register_fifo:fifo_data[0][6] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][6]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data06),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][6] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][6] .power_up = "low";

dffeas \register_fifo:fifo_data[0][7] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][7]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data07),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][7] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][7] .power_up = "low";

dffeas \register_fifo:fifo_data[0][8] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][8]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data08),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][8] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][8] .power_up = "low";

dffeas \register_fifo:fifo_data[0][9] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data09),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][9] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][9] .power_up = "low";

dffeas \register_fifo:fifo_data[0][10] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][10]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data010),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][10] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][10] .power_up = "low";

dffeas \register_fifo:fifo_data[0][11] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][11]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data011),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][11] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][11] .power_up = "low";

dffeas \register_fifo:fifo_data[0][12] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data012),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][12] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][12] .power_up = "low";

dffeas \register_fifo:fifo_data[0][13] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][13]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data013),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][13] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][13] .power_up = "low";

dffeas \register_fifo:fifo_data[0][14] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][14]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data014),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][14] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][14] .power_up = "low";

dffeas \register_fifo:fifo_data[0][15] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][15]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data015),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][15] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][15] .power_up = "low";

dffeas \register_fifo:fifo_data[0][16] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][16]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data016),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][16] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][16] .power_up = "low";

dffeas \register_fifo:fifo_data[0][17] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][17]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data017),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][17] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][17] .power_up = "low";

dffeas \register_fifo:fifo_data[0][18] (
	.clk(clk),
	.d(\register_fifo:fifo_data[0][18]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!enable),
	.q(register_fifofifo_data018),
	.prn(vcc));
defparam \register_fifo:fifo_data[0][18] .is_wysiwyg = "true";
defparam \register_fifo:fifo_data[0][18] .power_up = "low";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][0]~1 (
	.dataa(register_fifofifo_data00),
	.datab(register_fifofifo_data001),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\register_fifo:fifo_data[0][0]~1_combout ),
	.cout(\register_fifo:fifo_data[0][0]~2 ));
defparam \register_fifo:fifo_data[0][0]~1 .lut_mask = 16'h66EE;
defparam \register_fifo:fifo_data[0][0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][1]~1 (
	.dataa(register_fifofifo_data01),
	.datab(register_fifofifo_data019),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][0]~2 ),
	.combout(\register_fifo:fifo_data[0][1]~1_combout ),
	.cout(\register_fifo:fifo_data[0][1]~2 ));
defparam \register_fifo:fifo_data[0][1]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][1]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][2]~1 (
	.dataa(register_fifofifo_data02),
	.datab(register_fifofifo_data021),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][1]~2 ),
	.combout(\register_fifo:fifo_data[0][2]~1_combout ),
	.cout(\register_fifo:fifo_data[0][2]~2 ));
defparam \register_fifo:fifo_data[0][2]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][2]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][3]~1 (
	.dataa(register_fifofifo_data03),
	.datab(register_fifofifo_data031),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][2]~2 ),
	.combout(\register_fifo:fifo_data[0][3]~1_combout ),
	.cout(\register_fifo:fifo_data[0][3]~2 ));
defparam \register_fifo:fifo_data[0][3]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][3]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][4]~1 (
	.dataa(register_fifofifo_data04),
	.datab(register_fifofifo_data041),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][3]~2 ),
	.combout(\register_fifo:fifo_data[0][4]~1_combout ),
	.cout(\register_fifo:fifo_data[0][4]~2 ));
defparam \register_fifo:fifo_data[0][4]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][4]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][5]~1 (
	.dataa(register_fifofifo_data05),
	.datab(register_fifofifo_data051),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][4]~2 ),
	.combout(\register_fifo:fifo_data[0][5]~1_combout ),
	.cout(\register_fifo:fifo_data[0][5]~2 ));
defparam \register_fifo:fifo_data[0][5]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][5]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][6]~1 (
	.dataa(register_fifofifo_data06),
	.datab(register_fifofifo_data061),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][5]~2 ),
	.combout(\register_fifo:fifo_data[0][6]~1_combout ),
	.cout(\register_fifo:fifo_data[0][6]~2 ));
defparam \register_fifo:fifo_data[0][6]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][6]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][7]~1 (
	.dataa(register_fifofifo_data07),
	.datab(register_fifofifo_data071),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][6]~2 ),
	.combout(\register_fifo:fifo_data[0][7]~1_combout ),
	.cout(\register_fifo:fifo_data[0][7]~2 ));
defparam \register_fifo:fifo_data[0][7]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][7]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][8]~1 (
	.dataa(register_fifofifo_data08),
	.datab(register_fifofifo_data081),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][7]~2 ),
	.combout(\register_fifo:fifo_data[0][8]~1_combout ),
	.cout(\register_fifo:fifo_data[0][8]~2 ));
defparam \register_fifo:fifo_data[0][8]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][8]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][9]~1 (
	.dataa(register_fifofifo_data09),
	.datab(register_fifofifo_data091),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][8]~2 ),
	.combout(\register_fifo:fifo_data[0][9]~1_combout ),
	.cout(\register_fifo:fifo_data[0][9]~2 ));
defparam \register_fifo:fifo_data[0][9]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][9]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][10]~1 (
	.dataa(register_fifofifo_data010),
	.datab(register_fifofifo_data0101),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][9]~2 ),
	.combout(\register_fifo:fifo_data[0][10]~1_combout ),
	.cout(\register_fifo:fifo_data[0][10]~2 ));
defparam \register_fifo:fifo_data[0][10]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][10]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][11]~1 (
	.dataa(register_fifofifo_data011),
	.datab(register_fifofifo_data0111),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][10]~2 ),
	.combout(\register_fifo:fifo_data[0][11]~1_combout ),
	.cout(\register_fifo:fifo_data[0][11]~2 ));
defparam \register_fifo:fifo_data[0][11]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][11]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][12]~1 (
	.dataa(register_fifofifo_data012),
	.datab(register_fifofifo_data0121),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][11]~2 ),
	.combout(\register_fifo:fifo_data[0][12]~1_combout ),
	.cout(\register_fifo:fifo_data[0][12]~2 ));
defparam \register_fifo:fifo_data[0][12]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][12]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][13]~1 (
	.dataa(register_fifofifo_data013),
	.datab(register_fifofifo_data0131),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][12]~2 ),
	.combout(\register_fifo:fifo_data[0][13]~1_combout ),
	.cout(\register_fifo:fifo_data[0][13]~2 ));
defparam \register_fifo:fifo_data[0][13]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][13]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][14]~1 (
	.dataa(register_fifofifo_data014),
	.datab(register_fifofifo_data0141),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][13]~2 ),
	.combout(\register_fifo:fifo_data[0][14]~1_combout ),
	.cout(\register_fifo:fifo_data[0][14]~2 ));
defparam \register_fifo:fifo_data[0][14]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][14]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][15]~1 (
	.dataa(register_fifofifo_data015),
	.datab(register_fifofifo_data0151),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][14]~2 ),
	.combout(\register_fifo:fifo_data[0][15]~1_combout ),
	.cout(\register_fifo:fifo_data[0][15]~2 ));
defparam \register_fifo:fifo_data[0][15]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][15]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][16]~1 (
	.dataa(register_fifofifo_data016),
	.datab(register_fifofifo_data0161),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][15]~2 ),
	.combout(\register_fifo:fifo_data[0][16]~1_combout ),
	.cout(\register_fifo:fifo_data[0][16]~2 ));
defparam \register_fifo:fifo_data[0][16]~1 .lut_mask = 16'h96EF;
defparam \register_fifo:fifo_data[0][16]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][17]~1 (
	.dataa(register_fifofifo_data017),
	.datab(register_fifofifo_data0171),
	.datac(gnd),
	.datad(vcc),
	.cin(\register_fifo:fifo_data[0][16]~2 ),
	.combout(\register_fifo:fifo_data[0][17]~1_combout ),
	.cout(\register_fifo:fifo_data[0][17]~2 ));
defparam \register_fifo:fifo_data[0][17]~1 .lut_mask = 16'h967F;
defparam \register_fifo:fifo_data[0][17]~1 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \register_fifo:fifo_data[0][18]~1 (
	.dataa(register_fifofifo_data018),
	.datab(register_fifofifo_data0181),
	.datac(gnd),
	.datad(gnd),
	.cin(\register_fifo:fifo_data[0][17]~2 ),
	.combout(\register_fifo:fifo_data[0][18]~1_combout ),
	.cout());
defparam \register_fifo:fifo_data[0][18]~1 .lut_mask = 16'h9696;
defparam \register_fifo:fifo_data[0][18]~1 .sum_lutc_input = "cin";

endmodule

module cic_counter_module_19 (
	ena_sample,
	stall_reg,
	count_0,
	count_3,
	count_2,
	count_1,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	ena_sample;
input 	stall_reg;
output 	count_0;
output 	count_3;
output 	count_2;
output 	count_1;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \count[0]~0_combout ;
wire \count~1_combout ;
wire \count[0]~2_combout ;
wire \Add0~0_combout ;
wire \count~3_combout ;
wire \Add0~1_combout ;
wire \count~4_combout ;
wire \count~5_combout ;


dffeas \count[0] (
	.clk(clk),
	.d(\count~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count[0]~2_combout ),
	.q(count_0),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

dffeas \count[3] (
	.clk(clk),
	.d(\count~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count[0]~2_combout ),
	.q(count_3),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

dffeas \count[2] (
	.clk(clk),
	.d(\count~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count[0]~2_combout ),
	.q(count_2),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

dffeas \count[1] (
	.clk(clk),
	.d(\count~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\count[0]~2_combout ),
	.q(count_1),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

fiftyfivenm_lcell_comb \count[0]~0 (
	.dataa(count_1),
	.datab(count_2),
	.datac(count_0),
	.datad(count_3),
	.cin(gnd),
	.combout(\count[0]~0_combout ),
	.cout());
defparam \count[0]~0 .lut_mask = 16'hFEFF;
defparam \count[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \count~1 (
	.dataa(count_0),
	.datab(gnd),
	.datac(reset_n),
	.datad(\count[0]~0_combout ),
	.cin(gnd),
	.combout(\count~1_combout ),
	.cout());
defparam \count~1 .lut_mask = 16'hFFF5;
defparam \count~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \count[0]~2 (
	.dataa(reset_n),
	.datab(stall_reg),
	.datac(gnd),
	.datad(ena_sample),
	.cin(gnd),
	.combout(\count[0]~2_combout ),
	.cout());
defparam \count[0]~2 .lut_mask = 16'hFF77;
defparam \count[0]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~0 (
	.dataa(count_3),
	.datab(count_1),
	.datac(count_2),
	.datad(count_0),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
defparam \Add0~0 .lut_mask = 16'h6996;
defparam \Add0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \count~3 (
	.dataa(reset_n),
	.datab(\count[0]~0_combout ),
	.datac(\Add0~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~3_combout ),
	.cout());
defparam \count~3 .lut_mask = 16'hFEFE;
defparam \count~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(count_2),
	.datac(count_1),
	.datad(count_0),
	.cin(gnd),
	.combout(\Add0~1_combout ),
	.cout());
defparam \Add0~1 .lut_mask = 16'hC33C;
defparam \Add0~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \count~4 (
	.dataa(reset_n),
	.datab(\count[0]~0_combout ),
	.datac(\Add0~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\count~4_combout ),
	.cout());
defparam \count~4 .lut_mask = 16'hFEFE;
defparam \count~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \count~5 (
	.dataa(reset_n),
	.datab(\count[0]~0_combout ),
	.datac(count_1),
	.datad(count_0),
	.cin(gnd),
	.combout(\count~5_combout ),
	.cout());
defparam \count~5 .lut_mask = 16'hEFFE;
defparam \count~5 .sum_lutc_input = "datac";

endmodule

module cic_auk_dspip_avalon_streaming_controller (
	dffe_nae,
	dffe_af,
	usedw_process,
	sink_ready_ctrl,
	sink_ready_ctrl1,
	stall_reg1,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	dffe_nae;
input 	dffe_af;
output 	usedw_process;
output 	sink_ready_ctrl;
output 	sink_ready_ctrl1;
output 	stall_reg1;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ready_FIFO|fifo_array[5][0]~q ;
wire \ready_FIFO|fifo_array[4][0]~q ;
wire \ready_FIFO|rd_addr_ptr[2]~q ;
wire \ready_FIFO|rd_addr_ptr[0]~q ;
wire \ready_FIFO|rd_addr_ptr[1]~q ;
wire \ready_FIFO|Equal2~0_combout ;
wire \ready_FIFO|Mux0~1_combout ;
wire \sink_ready_ctrl~0_combout ;
wire \stall_reg~0_combout ;


cic_auk_dspip_avalon_streaming_small_fifo ready_FIFO(
	.dffe_nae(dffe_nae),
	.dffe_af(dffe_af),
	.fifo_array_0_5(\ready_FIFO|fifo_array[5][0]~q ),
	.fifo_array_0_4(\ready_FIFO|fifo_array[4][0]~q ),
	.rd_addr_ptr_2(\ready_FIFO|rd_addr_ptr[2]~q ),
	.usedw_process(usedw_process),
	.rd_addr_ptr_0(\ready_FIFO|rd_addr_ptr[0]~q ),
	.rd_addr_ptr_1(\ready_FIFO|rd_addr_ptr[1]~q ),
	.Equal2(\ready_FIFO|Equal2~0_combout ),
	.Mux0(\ready_FIFO|Mux0~1_combout ),
	.stall_reg(stall_reg1),
	.clock(clk),
	.reset_n(reset_n));

fiftyfivenm_lcell_comb \sink_ready_ctrl~1 (
	.dataa(\sink_ready_ctrl~0_combout ),
	.datab(\ready_FIFO|rd_addr_ptr[2]~q ),
	.datac(gnd),
	.datad(\ready_FIFO|rd_addr_ptr[1]~q ),
	.cin(gnd),
	.combout(sink_ready_ctrl),
	.cout());
defparam \sink_ready_ctrl~1 .lut_mask = 16'hEEFF;
defparam \sink_ready_ctrl~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \sink_ready_ctrl~2 (
	.dataa(\ready_FIFO|Equal2~0_combout ),
	.datab(\ready_FIFO|Mux0~1_combout ),
	.datac(gnd),
	.datad(\ready_FIFO|rd_addr_ptr[2]~q ),
	.cin(gnd),
	.combout(sink_ready_ctrl1),
	.cout());
defparam \sink_ready_ctrl~2 .lut_mask = 16'hEEFF;
defparam \sink_ready_ctrl~2 .sum_lutc_input = "datac";

dffeas stall_reg(
	.clk(clk),
	.d(\stall_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stall_reg1),
	.prn(vcc));
defparam stall_reg.is_wysiwyg = "true";
defparam stall_reg.power_up = "low";

fiftyfivenm_lcell_comb \sink_ready_ctrl~0 (
	.dataa(\ready_FIFO|fifo_array[5][0]~q ),
	.datab(\ready_FIFO|fifo_array[4][0]~q ),
	.datac(gnd),
	.datad(\ready_FIFO|rd_addr_ptr[0]~q ),
	.cin(gnd),
	.combout(\sink_ready_ctrl~0_combout ),
	.cout());
defparam \sink_ready_ctrl~0 .lut_mask = 16'hAACC;
defparam \sink_ready_ctrl~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \stall_reg~0 (
	.dataa(dffe_af),
	.datab(gnd),
	.datac(dffe_nae),
	.datad(reset_n),
	.cin(gnd),
	.combout(\stall_reg~0_combout ),
	.cout());
defparam \stall_reg~0 .lut_mask = 16'hAFFF;
defparam \stall_reg~0 .sum_lutc_input = "datac";

endmodule

module cic_auk_dspip_avalon_streaming_small_fifo (
	dffe_nae,
	dffe_af,
	fifo_array_0_5,
	fifo_array_0_4,
	rd_addr_ptr_2,
	usedw_process,
	rd_addr_ptr_0,
	rd_addr_ptr_1,
	Equal2,
	Mux0,
	stall_reg,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	dffe_nae;
input 	dffe_af;
output 	fifo_array_0_5;
output 	fifo_array_0_4;
output 	rd_addr_ptr_2;
output 	usedw_process;
output 	rd_addr_ptr_0;
output 	rd_addr_ptr_1;
output 	Equal2;
output 	Mux0;
input 	stall_reg;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_addr_ptr~2_combout ;
wire \fifo_usedw[2]~0_combout ;
wire \fifo_usedw[0]~2_combout ;
wire \fifo_usedw[0]~3_combout ;
wire \fifo_usedw[0]~q ;
wire \usedw_process~4_combout ;
wire \Add2~1_combout ;
wire \fifo_usedw[1]~4_combout ;
wire \fifo_usedw[1]~q ;
wire \Add2~0_combout ;
wire \fifo_usedw[2]~1_combout ;
wire \fifo_usedw[2]~q ;
wire \usedw_process~3_combout ;
wire \wr_addr_ptr[2]~1_combout ;
wire \wr_addr_ptr[0]~q ;
wire \wr_addr_ptr~3_combout ;
wire \wr_addr_ptr[2]~q ;
wire \wr_addr_ptr~0_combout ;
wire \wr_addr_ptr[1]~q ;
wire \Decoder0~0_combout ;
wire \fifo_array~0_combout ;
wire \fifo_array~1_combout ;
wire \rd_addr_ptr~3_combout ;
wire \rd_addr_ptr[0]~5_combout ;
wire \rd_addr_ptr~2_combout ;
wire \rd_addr_ptr~4_combout ;
wire \Decoder0~1_combout ;
wire \Decoder0~2_combout ;
wire \fifo_array~2_combout ;
wire \fifo_array[2][0]~q ;
wire \fifo_array~3_combout ;
wire \fifo_array[1][0]~q ;
wire \fifo_array~4_combout ;
wire \fifo_array[0][0]~q ;
wire \Mux0~0_combout ;
wire \fifo_array~5_combout ;
wire \fifo_array[3][0]~q ;


dffeas \fifo_array[5][0] (
	.clk(clock),
	.d(\fifo_array~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_array_0_5),
	.prn(vcc));
defparam \fifo_array[5][0] .is_wysiwyg = "true";
defparam \fifo_array[5][0] .power_up = "low";

dffeas \fifo_array[4][0] (
	.clk(clock),
	.d(\fifo_array~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(fifo_array_0_4),
	.prn(vcc));
defparam \fifo_array[4][0] .is_wysiwyg = "true";
defparam \fifo_array[4][0] .power_up = "low";

dffeas \rd_addr_ptr[2] (
	.clk(clock),
	.d(\rd_addr_ptr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\rd_addr_ptr[0]~5_combout ),
	.q(rd_addr_ptr_2),
	.prn(vcc));
defparam \rd_addr_ptr[2] .is_wysiwyg = "true";
defparam \rd_addr_ptr[2] .power_up = "low";

fiftyfivenm_lcell_comb \usedw_process~2 (
	.dataa(dffe_nae),
	.datab(gnd),
	.datac(gnd),
	.datad(dffe_af),
	.cin(gnd),
	.combout(usedw_process),
	.cout());
defparam \usedw_process~2 .lut_mask = 16'hAAFF;
defparam \usedw_process~2 .sum_lutc_input = "datac";

dffeas \rd_addr_ptr[0] (
	.clk(clock),
	.d(\rd_addr_ptr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_addr_ptr[0]~5_combout ),
	.q(rd_addr_ptr_0),
	.prn(vcc));
defparam \rd_addr_ptr[0] .is_wysiwyg = "true";
defparam \rd_addr_ptr[0] .power_up = "low";

dffeas \rd_addr_ptr[1] (
	.clk(clock),
	.d(\rd_addr_ptr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_addr_ptr[0]~5_combout ),
	.q(rd_addr_ptr_1),
	.prn(vcc));
defparam \rd_addr_ptr[1] .is_wysiwyg = "true";
defparam \rd_addr_ptr[1] .power_up = "low";

fiftyfivenm_lcell_comb \Equal2~0 (
	.dataa(gnd),
	.datab(\fifo_usedw[2]~q ),
	.datac(\fifo_usedw[0]~q ),
	.datad(\fifo_usedw[1]~q ),
	.cin(gnd),
	.combout(Equal2),
	.cout());
defparam \Equal2~0 .lut_mask = 16'h3FFF;
defparam \Equal2~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Mux0~1 (
	.dataa(\fifo_array[2][0]~q ),
	.datab(rd_addr_ptr_1),
	.datac(\Mux0~0_combout ),
	.datad(\fifo_array[3][0]~q ),
	.cin(gnd),
	.combout(Mux0),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hFFBE;
defparam \Mux0~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \wr_addr_ptr~2 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\wr_addr_ptr[0]~q ),
	.cin(gnd),
	.combout(\wr_addr_ptr~2_combout ),
	.cout());
defparam \wr_addr_ptr~2 .lut_mask = 16'hAAFF;
defparam \wr_addr_ptr~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \fifo_usedw[2]~0 (
	.dataa(usedw_process),
	.datab(\usedw_process~3_combout ),
	.datac(Equal2),
	.datad(reset_n),
	.cin(gnd),
	.combout(\fifo_usedw[2]~0_combout ),
	.cout());
defparam \fifo_usedw[2]~0 .lut_mask = 16'h6FFF;
defparam \fifo_usedw[2]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \fifo_usedw[0]~2 (
	.dataa(\fifo_usedw[0]~q ),
	.datab(Equal2),
	.datac(usedw_process),
	.datad(\usedw_process~3_combout ),
	.cin(gnd),
	.combout(\fifo_usedw[0]~2_combout ),
	.cout());
defparam \fifo_usedw[0]~2 .lut_mask = 16'h6996;
defparam \fifo_usedw[0]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \fifo_usedw[0]~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(reset_n),
	.datad(\fifo_usedw[0]~2_combout ),
	.cin(gnd),
	.combout(\fifo_usedw[0]~3_combout ),
	.cout());
defparam \fifo_usedw[0]~3 .lut_mask = 16'hFFF0;
defparam \fifo_usedw[0]~3 .sum_lutc_input = "datac";

dffeas \fifo_usedw[0] (
	.clk(clock),
	.d(\fifo_usedw[0]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_usedw[0]~q ),
	.prn(vcc));
defparam \fifo_usedw[0] .is_wysiwyg = "true";
defparam \fifo_usedw[0] .power_up = "low";

fiftyfivenm_lcell_comb \usedw_process~4 (
	.dataa(dffe_nae),
	.datab(dffe_af),
	.datac(\usedw_process~3_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\usedw_process~4_combout ),
	.cout());
defparam \usedw_process~4 .lut_mask = 16'hDFDF;
defparam \usedw_process~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add2~1 (
	.dataa(\fifo_usedw[0]~q ),
	.datab(\fifo_usedw[1]~q ),
	.datac(\usedw_process~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add2~1_combout ),
	.cout());
defparam \Add2~1 .lut_mask = 16'h9696;
defparam \Add2~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \fifo_usedw[1]~4 (
	.dataa(\fifo_usedw[1]~q ),
	.datab(reset_n),
	.datac(\fifo_usedw[2]~0_combout ),
	.datad(\Add2~1_combout ),
	.cin(gnd),
	.combout(\fifo_usedw[1]~4_combout ),
	.cout());
defparam \fifo_usedw[1]~4 .lut_mask = 16'hACFF;
defparam \fifo_usedw[1]~4 .sum_lutc_input = "datac";

dffeas \fifo_usedw[1] (
	.clk(clock),
	.d(\fifo_usedw[1]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_usedw[1]~q ),
	.prn(vcc));
defparam \fifo_usedw[1] .is_wysiwyg = "true";
defparam \fifo_usedw[1] .power_up = "low";

fiftyfivenm_lcell_comb \Add2~0 (
	.dataa(\fifo_usedw[0]~q ),
	.datab(\fifo_usedw[1]~q ),
	.datac(\usedw_process~4_combout ),
	.datad(\fifo_usedw[2]~q ),
	.cin(gnd),
	.combout(\Add2~0_combout ),
	.cout());
defparam \Add2~0 .lut_mask = 16'h6996;
defparam \Add2~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \fifo_usedw[2]~1 (
	.dataa(\fifo_usedw[2]~q ),
	.datab(reset_n),
	.datac(\fifo_usedw[2]~0_combout ),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\fifo_usedw[2]~1_combout ),
	.cout());
defparam \fifo_usedw[2]~1 .lut_mask = 16'hACFF;
defparam \fifo_usedw[2]~1 .sum_lutc_input = "datac";

dffeas \fifo_usedw[2] (
	.clk(clock),
	.d(\fifo_usedw[2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_usedw[2]~q ),
	.prn(vcc));
defparam \fifo_usedw[2] .is_wysiwyg = "true";
defparam \fifo_usedw[2] .power_up = "low";

fiftyfivenm_lcell_comb \usedw_process~3 (
	.dataa(stall_reg),
	.datab(\fifo_usedw[2]~q ),
	.datac(\fifo_usedw[1]~q ),
	.datad(\fifo_usedw[0]~q ),
	.cin(gnd),
	.combout(\usedw_process~3_combout ),
	.cout());
defparam \usedw_process~3 .lut_mask = 16'hFEFF;
defparam \usedw_process~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \wr_addr_ptr[2]~1 (
	.dataa(reset_n),
	.datab(\usedw_process~3_combout ),
	.datac(usedw_process),
	.datad(Equal2),
	.cin(gnd),
	.combout(\wr_addr_ptr[2]~1_combout ),
	.cout());
defparam \wr_addr_ptr[2]~1 .lut_mask = 16'h7FFF;
defparam \wr_addr_ptr[2]~1 .sum_lutc_input = "datac";

dffeas \wr_addr_ptr[0] (
	.clk(clock),
	.d(\wr_addr_ptr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_addr_ptr[2]~1_combout ),
	.q(\wr_addr_ptr[0]~q ),
	.prn(vcc));
defparam \wr_addr_ptr[0] .is_wysiwyg = "true";
defparam \wr_addr_ptr[0] .power_up = "low";

fiftyfivenm_lcell_comb \wr_addr_ptr~3 (
	.dataa(\wr_addr_ptr[1]~q ),
	.datab(gnd),
	.datac(\wr_addr_ptr[2]~q ),
	.datad(\wr_addr_ptr[0]~q ),
	.cin(gnd),
	.combout(\wr_addr_ptr~3_combout ),
	.cout());
defparam \wr_addr_ptr~3 .lut_mask = 16'hAFFA;
defparam \wr_addr_ptr~3 .sum_lutc_input = "datac";

dffeas \wr_addr_ptr[2] (
	.clk(clock),
	.d(\wr_addr_ptr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(\wr_addr_ptr[2]~1_combout ),
	.q(\wr_addr_ptr[2]~q ),
	.prn(vcc));
defparam \wr_addr_ptr[2] .is_wysiwyg = "true";
defparam \wr_addr_ptr[2] .power_up = "low";

fiftyfivenm_lcell_comb \wr_addr_ptr~0 (
	.dataa(reset_n),
	.datab(\wr_addr_ptr[1]~q ),
	.datac(\wr_addr_ptr[2]~q ),
	.datad(\wr_addr_ptr[0]~q ),
	.cin(gnd),
	.combout(\wr_addr_ptr~0_combout ),
	.cout());
defparam \wr_addr_ptr~0 .lut_mask = 16'hBFEF;
defparam \wr_addr_ptr~0 .sum_lutc_input = "datac";

dffeas \wr_addr_ptr[1] (
	.clk(clock),
	.d(\wr_addr_ptr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_addr_ptr[2]~1_combout ),
	.q(\wr_addr_ptr[1]~q ),
	.prn(vcc));
defparam \wr_addr_ptr[1] .is_wysiwyg = "true";
defparam \wr_addr_ptr[1] .power_up = "low";

fiftyfivenm_lcell_comb \Decoder0~0 (
	.dataa(usedw_process),
	.datab(Equal2),
	.datac(\wr_addr_ptr[1]~q ),
	.datad(\usedw_process~3_combout ),
	.cin(gnd),
	.combout(\Decoder0~0_combout ),
	.cout());
defparam \Decoder0~0 .lut_mask = 16'h7FFF;
defparam \Decoder0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \fifo_array~0 (
	.dataa(fifo_array_0_5),
	.datab(\Decoder0~0_combout ),
	.datac(\wr_addr_ptr[0]~q ),
	.datad(\wr_addr_ptr[2]~q ),
	.cin(gnd),
	.combout(\fifo_array~0_combout ),
	.cout());
defparam \fifo_array~0 .lut_mask = 16'hFFFE;
defparam \fifo_array~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \fifo_array~1 (
	.dataa(fifo_array_0_4),
	.datab(\Decoder0~0_combout ),
	.datac(\wr_addr_ptr[2]~q ),
	.datad(\wr_addr_ptr[0]~q ),
	.cin(gnd),
	.combout(\fifo_array~1_combout ),
	.cout());
defparam \fifo_array~1 .lut_mask = 16'hFEFF;
defparam \fifo_array~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_addr_ptr~3 (
	.dataa(rd_addr_ptr_1),
	.datab(gnd),
	.datac(rd_addr_ptr_2),
	.datad(rd_addr_ptr_0),
	.cin(gnd),
	.combout(\rd_addr_ptr~3_combout ),
	.cout());
defparam \rd_addr_ptr~3 .lut_mask = 16'hAFFA;
defparam \rd_addr_ptr~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_addr_ptr[0]~5 (
	.dataa(dffe_nae),
	.datab(dffe_af),
	.datac(reset_n),
	.datad(Equal2),
	.cin(gnd),
	.combout(\rd_addr_ptr[0]~5_combout ),
	.cout());
defparam \rd_addr_ptr[0]~5 .lut_mask = 16'hBFFF;
defparam \rd_addr_ptr[0]~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_addr_ptr~2 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(rd_addr_ptr_0),
	.cin(gnd),
	.combout(\rd_addr_ptr~2_combout ),
	.cout());
defparam \rd_addr_ptr~2 .lut_mask = 16'hAAFF;
defparam \rd_addr_ptr~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_addr_ptr~4 (
	.dataa(reset_n),
	.datab(rd_addr_ptr_1),
	.datac(rd_addr_ptr_2),
	.datad(rd_addr_ptr_0),
	.cin(gnd),
	.combout(\rd_addr_ptr~4_combout ),
	.cout());
defparam \rd_addr_ptr~4 .lut_mask = 16'hBFEF;
defparam \rd_addr_ptr~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Decoder0~1 (
	.dataa(\wr_addr_ptr[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\wr_addr_ptr[2]~q ),
	.cin(gnd),
	.combout(\Decoder0~1_combout ),
	.cout());
defparam \Decoder0~1 .lut_mask = 16'hAAFF;
defparam \Decoder0~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Decoder0~2 (
	.dataa(\Decoder0~1_combout ),
	.datab(usedw_process),
	.datac(Equal2),
	.datad(\usedw_process~3_combout ),
	.cin(gnd),
	.combout(\Decoder0~2_combout ),
	.cout());
defparam \Decoder0~2 .lut_mask = 16'hBFFF;
defparam \Decoder0~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \fifo_array~2 (
	.dataa(\fifo_array[2][0]~q ),
	.datab(\Decoder0~2_combout ),
	.datac(gnd),
	.datad(\wr_addr_ptr[0]~q ),
	.cin(gnd),
	.combout(\fifo_array~2_combout ),
	.cout());
defparam \fifo_array~2 .lut_mask = 16'hEEFF;
defparam \fifo_array~2 .sum_lutc_input = "datac";

dffeas \fifo_array[2][0] (
	.clk(clock),
	.d(\fifo_array~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_array[2][0]~q ),
	.prn(vcc));
defparam \fifo_array[2][0] .is_wysiwyg = "true";
defparam \fifo_array[2][0] .power_up = "low";

fiftyfivenm_lcell_comb \fifo_array~3 (
	.dataa(\fifo_array[1][0]~q ),
	.datab(\Decoder0~0_combout ),
	.datac(\wr_addr_ptr[0]~q ),
	.datad(\wr_addr_ptr[2]~q ),
	.cin(gnd),
	.combout(\fifo_array~3_combout ),
	.cout());
defparam \fifo_array~3 .lut_mask = 16'hFEFF;
defparam \fifo_array~3 .sum_lutc_input = "datac";

dffeas \fifo_array[1][0] (
	.clk(clock),
	.d(\fifo_array~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_array[1][0]~q ),
	.prn(vcc));
defparam \fifo_array[1][0] .is_wysiwyg = "true";
defparam \fifo_array[1][0] .power_up = "low";

fiftyfivenm_lcell_comb \fifo_array~4 (
	.dataa(\fifo_array[0][0]~q ),
	.datab(\Decoder0~0_combout ),
	.datac(\wr_addr_ptr[0]~q ),
	.datad(\wr_addr_ptr[2]~q ),
	.cin(gnd),
	.combout(\fifo_array~4_combout ),
	.cout());
defparam \fifo_array~4 .lut_mask = 16'hEFFF;
defparam \fifo_array~4 .sum_lutc_input = "datac";

dffeas \fifo_array[0][0] (
	.clk(clock),
	.d(\fifo_array~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_array[0][0]~q ),
	.prn(vcc));
defparam \fifo_array[0][0] .is_wysiwyg = "true";
defparam \fifo_array[0][0] .power_up = "low";

fiftyfivenm_lcell_comb \Mux0~0 (
	.dataa(rd_addr_ptr_1),
	.datab(\fifo_array[1][0]~q ),
	.datac(rd_addr_ptr_0),
	.datad(\fifo_array[0][0]~q ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hFFDE;
defparam \Mux0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \fifo_array~5 (
	.dataa(\fifo_array[3][0]~q ),
	.datab(\wr_addr_ptr[0]~q ),
	.datac(\Decoder0~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_array~5_combout ),
	.cout());
defparam \fifo_array~5 .lut_mask = 16'hFEFE;
defparam \fifo_array~5 .sum_lutc_input = "datac";

dffeas \fifo_array[3][0] (
	.clk(clock),
	.d(\fifo_array~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_array[3][0]~q ),
	.prn(vcc));
defparam \fifo_array[3][0] .is_wysiwyg = "true";
defparam \fifo_array[3][0] .power_up = "low";

endmodule

module cic_auk_dspip_avalon_streaming_sink (
	full_dff,
	dffe_nae,
	dffe_af,
	data,
	usedw_process,
	sink_ready_ctrl,
	sink_ready_ctrl1,
	GND_port,
	clk,
	in_valid,
	reset_n,
	at_sink_data)/* synthesis synthesis_greybox=1 */;
output 	full_dff;
output 	dffe_nae;
input 	dffe_af;
output 	[8:0] data;
input 	usedw_process;
input 	sink_ready_ctrl;
input 	sink_ready_ctrl1;
input 	GND_port;
input 	clk;
input 	in_valid;
input 	reset_n;
input 	[8:0] at_sink_data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_10 sink_FIFO(
	.full_dff(full_dff),
	.dffe_nae(dffe_nae),
	.dffe_af(dffe_af),
	.q({q_unconnected_wire_22,q_unconnected_wire_21,q_unconnected_wire_20,q_unconnected_wire_19,q_unconnected_wire_18,q_unconnected_wire_17,q_unconnected_wire_16,q_unconnected_wire_15,q_unconnected_wire_14,q_unconnected_wire_13,q_unconnected_wire_12,q_unconnected_wire_11,
q_unconnected_wire_10,q_unconnected_wire_9,data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.usedw_process(usedw_process),
	.sink_ready_ctrl(sink_ready_ctrl),
	.sink_ready_ctrl1(sink_ready_ctrl1),
	.GND_port(GND_port),
	.clock(clk),
	.in_valid(in_valid),
	.reset_n(reset_n),
	.data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,at_sink_data[8],at_sink_data[7],at_sink_data[6],at_sink_data[5],at_sink_data[4],at_sink_data[3],at_sink_data[2],at_sink_data[1],at_sink_data[0]}));

endmodule

module cic_scfifo_10 (
	full_dff,
	dffe_nae,
	dffe_af,
	q,
	usedw_process,
	sink_ready_ctrl,
	sink_ready_ctrl1,
	GND_port,
	clock,
	in_valid,
	reset_n,
	data)/* synthesis synthesis_greybox=1 */;
output 	full_dff;
output 	dffe_nae;
input 	dffe_af;
output 	[22:0] q;
input 	usedw_process;
input 	sink_ready_ctrl;
input 	sink_ready_ctrl1;
input 	GND_port;
input 	clock;
input 	in_valid;
input 	reset_n;
input 	[22:0] data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_vp61 auto_generated(
	.full_dff(full_dff),
	.dffe_nae1(dffe_nae),
	.dffe_af(dffe_af),
	.q({q_unconnected_wire_10,q_unconnected_wire_9,q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.usedw_process(usedw_process),
	.sink_ready_ctrl(sink_ready_ctrl),
	.sink_ready_ctrl1(sink_ready_ctrl1),
	.GND_port(GND_port),
	.clock(clock),
	.in_valid(in_valid),
	.reset_n(reset_n),
	.data({gnd,gnd,data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}));

endmodule

module cic_scfifo_vp61 (
	full_dff,
	dffe_nae1,
	dffe_af,
	q,
	usedw_process,
	sink_ready_ctrl,
	sink_ready_ctrl1,
	GND_port,
	clock,
	in_valid,
	reset_n,
	data)/* synthesis synthesis_greybox=1 */;
output 	full_dff;
output 	dffe_nae1;
input 	dffe_af;
output 	[10:0] q;
input 	usedw_process;
input 	sink_ready_ctrl;
input 	sink_ready_ctrl1;
input 	GND_port;
input 	clock;
input 	in_valid;
input 	reset_n;
input 	[10:0] data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dpfifo|usedw_counter|counter_reg_bit[2]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[1]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[0]~q ;
wire \dffe_nae~0_combout ;
wire \dffe_nae~1_combout ;
wire \dffe_nae~2_combout ;


cic_a_dpfifo_gvu dpfifo(
	.full_dff1(full_dff),
	.counter_reg_bit_2(\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.q({q_unconnected_wire_10,q_unconnected_wire_9,q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.usedw_process(usedw_process),
	.sink_ready_ctrl(sink_ready_ctrl),
	.sink_ready_ctrl1(sink_ready_ctrl1),
	.GND_port(GND_port),
	.clock(clock),
	.in_valid(in_valid),
	.reset_n(reset_n),
	.data({gnd,gnd,data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}));

dffeas dffe_nae(
	.clk(clock),
	.d(\dffe_nae~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(dffe_nae1),
	.prn(vcc));
defparam dffe_nae.is_wysiwyg = "true";
defparam dffe_nae.power_up = "low";

fiftyfivenm_lcell_comb \dffe_nae~0 (
	.dataa(sink_ready_ctrl),
	.datab(sink_ready_ctrl1),
	.datac(dffe_af),
	.datad(gnd),
	.cin(gnd),
	.combout(\dffe_nae~0_combout ),
	.cout());
defparam \dffe_nae~0 .lut_mask = 16'hEFEF;
defparam \dffe_nae~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dffe_nae~1 (
	.dataa(\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.datab(\dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.datac(\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.datad(dffe_nae1),
	.cin(gnd),
	.combout(\dffe_nae~1_combout ),
	.cout());
defparam \dffe_nae~1 .lut_mask = 16'h6996;
defparam \dffe_nae~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dffe_nae~2 (
	.dataa(in_valid),
	.datab(\dffe_nae~0_combout ),
	.datac(dffe_nae1),
	.datad(\dffe_nae~1_combout ),
	.cin(gnd),
	.combout(\dffe_nae~2_combout ),
	.cout());
defparam \dffe_nae~2 .lut_mask = 16'hBBF3;
defparam \dffe_nae~2 .sum_lutc_input = "datac";

endmodule

module cic_a_dpfifo_gvu (
	full_dff1,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	q,
	usedw_process,
	sink_ready_ctrl,
	sink_ready_ctrl1,
	GND_port,
	clock,
	in_valid,
	reset_n,
	data)/* synthesis synthesis_greybox=1 */;
output 	full_dff1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	[10:0] q;
input 	usedw_process;
input 	sink_ready_ctrl;
input 	sink_ready_ctrl1;
input 	GND_port;
input 	clock;
input 	in_valid;
input 	reset_n;
input 	[10:0] data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \_~0_combout ;
wire \empty_dff~2_combout ;
wire \usedw_is_0_dff~q ;
wire \valid_wreq~combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \empty_dff~1_combout ;
wire \empty_dff~q ;
wire \valid_rreq~combout ;
wire \_~1_combout ;


cic_cntr_hka rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.valid_rreq(\valid_rreq~combout ),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_altsyncram_thg1 FIFOram(
	.q_b({q_b_unconnected_wire_10,q_b_unconnected_wire_9,q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.address_a({\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.clocken1(\valid_rreq~combout ),
	.wren_a(\valid_wreq~combout ),
	.address_b({\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock0(clock),
	.clock1(clock),
	.data_a({gnd,gnd,data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}));

cic_cntr_ika_9 wr_ptr(
	.full_dff(full_dff1),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.GND_port(GND_port),
	.clock(clock),
	.in_valid(in_valid),
	.reset_n(reset_n));

cic_cntr_uk6 usedw_counter(
	.full_dff(full_dff1),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.valid_rreq(\valid_rreq~combout ),
	.updown(\valid_wreq~combout ),
	.GND_port(GND_port),
	.clock(clock),
	.in_valid(in_valid),
	.reset_n(reset_n));

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(\valid_rreq~combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(\valid_rreq~combout ),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(\valid_rreq~combout ),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(\valid_rreq~combout ),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~1 (
	.dataa(\valid_rreq~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(\valid_rreq~combout ),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(\valid_rreq~combout ),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

dffeas full_dff(
	.clk(clock),
	.d(\_~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(full_dff1),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(counter_reg_bit_2),
	.datab(in_valid),
	.datac(counter_reg_bit_1),
	.datad(counter_reg_bit_0),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hFFFE;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

fiftyfivenm_lcell_comb valid_wreq(
	.dataa(in_valid),
	.datab(gnd),
	.datac(gnd),
	.datad(full_dff1),
	.cin(gnd),
	.combout(\valid_wreq~combout ),
	.cout());
defparam valid_wreq.lut_mask = 16'hAAFF;
defparam valid_wreq.sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~0 (
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(counter_reg_bit_2),
	.datad(counter_reg_bit_0),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'hAFFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~1 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\valid_rreq~combout ),
	.datac(\usedw_will_be_1~0_combout ),
	.datad(\valid_wreq~combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFBFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~2 (
	.dataa(in_valid),
	.datab(gnd),
	.datac(full_dff1),
	.datad(\usedw_is_0_dff~q ),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hAFFF;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\usedw_will_be_1~2_combout ),
	.datad(\valid_rreq~combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFEFF;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

fiftyfivenm_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~combout ),
	.datac(\usedw_is_1_dff~q ),
	.datad(\valid_rreq~combout ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBFEF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hEFFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty_dff~q ),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

fiftyfivenm_lcell_comb valid_rreq(
	.dataa(\empty_dff~q ),
	.datab(usedw_process),
	.datac(sink_ready_ctrl),
	.datad(sink_ready_ctrl1),
	.cin(gnd),
	.combout(\valid_rreq~combout ),
	.cout());
defparam valid_rreq.lut_mask = 16'hFFFE;
defparam valid_rreq.sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \_~1 (
	.dataa(full_dff1),
	.datab(\_~0_combout ),
	.datac(gnd),
	.datad(\valid_rreq~combout ),
	.cin(gnd),
	.combout(\_~1_combout ),
	.cout());
defparam \_~1 .lut_mask = 16'hEEFF;
defparam \_~1 .sum_lutc_input = "datac";

endmodule

module cic_altsyncram_thg1 (
	q_b,
	address_a,
	clocken1,
	wren_a,
	address_b,
	clock0,
	clock1,
	data_a)/* synthesis synthesis_greybox=1 */;
output 	[10:0] q_b;
input 	[2:0] address_a;
input 	clocken1;
input 	wren_a;
input 	[2:0] address_b;
input 	clock0;
input 	clock1;
input 	[10:0] data_a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

fiftyfivenm_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_vp61:auto_generated|a_dpfifo_gvu:dpfifo|altsyncram_thg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 3;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 7;
defparam ram_block1a5.port_a_logical_ram_depth = 8;
defparam ram_block1a5.port_a_logical_ram_width = 11;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 3;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 7;
defparam ram_block1a5.port_b_logical_ram_depth = 8;
defparam ram_block1a5.port_b_logical_ram_width = 11;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_vp61:auto_generated|a_dpfifo_gvu:dpfifo|altsyncram_thg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 3;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 7;
defparam ram_block1a6.port_a_logical_ram_depth = 8;
defparam ram_block1a6.port_a_logical_ram_width = 11;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 3;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 7;
defparam ram_block1a6.port_b_logical_ram_depth = 8;
defparam ram_block1a6.port_b_logical_ram_width = 11;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk1_output_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_vp61:auto_generated|a_dpfifo_gvu:dpfifo|altsyncram_thg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 3;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 7;
defparam ram_block1a4.port_a_logical_ram_depth = 8;
defparam ram_block1a4.port_a_logical_ram_width = 11;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 3;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 7;
defparam ram_block1a4.port_b_logical_ram_depth = 8;
defparam ram_block1a4.port_b_logical_ram_width = 11;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_vp61:auto_generated|a_dpfifo_gvu:dpfifo|altsyncram_thg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 3;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 7;
defparam ram_block1a7.port_a_logical_ram_depth = 8;
defparam ram_block1a7.port_a_logical_ram_width = 11;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 3;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 7;
defparam ram_block1a7.port_b_logical_ram_depth = 8;
defparam ram_block1a7.port_b_logical_ram_width = 11;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk1_output_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_vp61:auto_generated|a_dpfifo_gvu:dpfifo|altsyncram_thg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 3;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 7;
defparam ram_block1a2.port_a_logical_ram_depth = 8;
defparam ram_block1a2.port_a_logical_ram_width = 11;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 3;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 7;
defparam ram_block1a2.port_b_logical_ram_depth = 8;
defparam ram_block1a2.port_b_logical_ram_width = 11;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk1_output_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_vp61:auto_generated|a_dpfifo_gvu:dpfifo|altsyncram_thg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 3;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 7;
defparam ram_block1a1.port_a_logical_ram_depth = 8;
defparam ram_block1a1.port_a_logical_ram_width = 11;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 3;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 7;
defparam ram_block1a1.port_b_logical_ram_depth = 8;
defparam ram_block1a1.port_b_logical_ram_width = 11;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk1_output_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_vp61:auto_generated|a_dpfifo_gvu:dpfifo|altsyncram_thg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 3;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 7;
defparam ram_block1a0.port_a_logical_ram_depth = 8;
defparam ram_block1a0.port_a_logical_ram_width = 11;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 3;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 7;
defparam ram_block1a0.port_b_logical_ram_depth = 8;
defparam ram_block1a0.port_b_logical_ram_width = 11;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk1_output_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_vp61:auto_generated|a_dpfifo_gvu:dpfifo|altsyncram_thg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 3;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 7;
defparam ram_block1a3.port_a_logical_ram_depth = 8;
defparam ram_block1a3.port_a_logical_ram_width = 11;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 3;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 7;
defparam ram_block1a3.port_b_logical_ram_depth = 8;
defparam ram_block1a3.port_b_logical_ram_width = 11;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_sink:input_sink|scfifo:sink_FIFO|scfifo_vp61:auto_generated|a_dpfifo_gvu:dpfifo|altsyncram_thg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 3;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 7;
defparam ram_block1a8.port_a_logical_ram_depth = 8;
defparam ram_block1a8.port_a_logical_ram_width = 11;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 3;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 7;
defparam ram_block1a8.port_b_logical_ram_depth = 8;
defparam ram_block1a8.port_b_logical_ram_width = 11;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

endmodule

module cic_cntr_hka (
	counter_reg_bit_0,
	counter_reg_bit_1,
	valid_rreq,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
input 	valid_rreq;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(valid_rreq),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout());
defparam counter_comb_bita1.lut_mask = 16'h5A5A;
defparam counter_comb_bita1.sum_lutc_input = "cin";

endmodule

module cic_cntr_ika_9 (
	full_dff,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	GND_port,
	clock,
	in_valid,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
input 	GND_port;
input 	clock;
input 	in_valid;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(in_valid),
	.datab(gnd),
	.datac(full_dff),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout());
defparam counter_comb_bita2.lut_mask = 16'h5A5A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

endmodule

module cic_cntr_uk6 (
	full_dff,
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	valid_rreq,
	updown,
	GND_port,
	clock,
	in_valid,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	full_dff;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
input 	valid_rreq;
input 	updown;
input 	GND_port;
input 	clock;
input 	in_valid;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \_~2_combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~2_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout());
defparam counter_comb_bita2.lut_mask = 16'h5A5A;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~2 (
	.dataa(in_valid),
	.datab(full_dff),
	.datac(valid_rreq),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'h96FF;
defparam \_~2 .sum_lutc_input = "datac";

endmodule

module cic_auk_dspip_avalon_streaming_source (
	at_source_data,
	source_valid_s1,
	at_source_channel,
	dffe_af,
	state_0,
	data,
	Equal0,
	Equal1,
	stall_reg,
	dout_valid,
	data_count,
	GND_port,
	clk,
	reset_n,
	out_ready)/* synthesis synthesis_greybox=1 */;
output 	[18:0] at_source_data;
output 	source_valid_s1;
output 	[3:0] at_source_channel;
output 	dffe_af;
input 	state_0;
input 	[18:0] data;
output 	Equal0;
output 	Equal1;
input 	stall_reg;
input 	dout_valid;
input 	[3:0] data_count;
input 	GND_port;
input 	clk;
input 	reset_n;
input 	out_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \source_FIFO|auto_generated|dpfifo|empty_dff~q ;
wire \source_valid_s_process~0_combout ;
wire \source_valid_s_process~1_combout ;


cic_scfifo_11 source_FIFO(
	.q({at_source_channel[3],at_source_channel[2],at_source_channel[1],at_source_channel[0],at_source_data[18],at_source_data[17],at_source_data[16],at_source_data[15],at_source_data[14],at_source_data[13],at_source_data[12],at_source_data[11],at_source_data[10],at_source_data[9],at_source_data[8],at_source_data[7],at_source_data[6],
at_source_data[5],at_source_data[4],at_source_data[3],at_source_data[2],at_source_data[1],at_source_data[0]}),
	.source_valid_s(source_valid_s1),
	.dffe_af(dffe_af),
	.state_0(state_0),
	.data({data_count[3],data_count[2],data_count[1],data_count[0],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.dout_valid(dout_valid),
	.empty_dff(\source_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.source_valid_s_process(\source_valid_s_process~0_combout ),
	.GND_port(GND_port),
	.clock(clk),
	.reset_n(reset_n),
	.out_ready(out_ready));

fiftyfivenm_lcell_comb \source_valid_s_process~0 (
	.dataa(\source_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.datab(out_ready),
	.datac(gnd),
	.datad(source_valid_s1),
	.cin(gnd),
	.combout(\source_valid_s_process~0_combout ),
	.cout());
defparam \source_valid_s_process~0 .lut_mask = 16'hEEFF;
defparam \source_valid_s_process~0 .sum_lutc_input = "datac";

dffeas source_valid_s(
	.clk(clk),
	.d(\source_valid_s_process~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(source_valid_s1),
	.prn(vcc));
defparam source_valid_s.is_wysiwyg = "true";
defparam source_valid_s.power_up = "low";

fiftyfivenm_lcell_comb \Equal0~0 (
	.dataa(at_source_channel[3]),
	.datab(at_source_channel[0]),
	.datac(at_source_channel[1]),
	.datad(at_source_channel[2]),
	.cin(gnd),
	.combout(Equal0),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h7FFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal1~0 (
	.dataa(at_source_channel[3]),
	.datab(at_source_channel[0]),
	.datac(at_source_channel[1]),
	.datad(at_source_channel[2]),
	.cin(gnd),
	.combout(Equal1),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hBFFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \source_valid_s_process~1 (
	.dataa(out_ready),
	.datab(gnd),
	.datac(source_valid_s1),
	.datad(\source_FIFO|auto_generated|dpfifo|empty_dff~q ),
	.cin(gnd),
	.combout(\source_valid_s_process~1_combout ),
	.cout());
defparam \source_valid_s_process~1 .lut_mask = 16'hFFF5;
defparam \source_valid_s_process~1 .sum_lutc_input = "datac";

endmodule

module cic_scfifo_11 (
	q,
	source_valid_s,
	dffe_af,
	state_0,
	data,
	stall_reg,
	dout_valid,
	empty_dff,
	source_valid_s_process,
	GND_port,
	clock,
	reset_n,
	out_ready)/* synthesis synthesis_greybox=1 */;
output 	[22:0] q;
input 	source_valid_s;
output 	dffe_af;
input 	state_0;
input 	[22:0] data;
input 	stall_reg;
input 	dout_valid;
output 	empty_dff;
input 	source_valid_s_process;
input 	GND_port;
input 	clock;
input 	reset_n;
input 	out_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cic_scfifo_vs61 auto_generated(
	.q({q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.source_valid_s(source_valid_s),
	.dffe_af1(dffe_af),
	.state_0(state_0),
	.data({data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.stall_reg(stall_reg),
	.dout_valid(dout_valid),
	.empty_dff(empty_dff),
	.source_valid_s_process(source_valid_s_process),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n),
	.out_ready(out_ready));

endmodule

module cic_scfifo_vs61 (
	q,
	source_valid_s,
	dffe_af1,
	state_0,
	data,
	stall_reg,
	dout_valid,
	empty_dff,
	source_valid_s_process,
	GND_port,
	clock,
	reset_n,
	out_ready)/* synthesis synthesis_greybox=1 */;
output 	[22:0] q;
input 	source_valid_s;
output 	dffe_af1;
input 	state_0;
input 	[22:0] data;
input 	stall_reg;
input 	dout_valid;
output 	empty_dff;
input 	source_valid_s_process;
input 	GND_port;
input 	clock;
input 	reset_n;
input 	out_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dpfifo|usedw_counter|counter_reg_bit[2]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[3]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[1]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[4]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[0]~q ;
wire \dffe_af~0_combout ;
wire \dffe_af~1_combout ;
wire \dffe_af~2_combout ;
wire \dffe_af~3_combout ;


cic_a_dpfifo_s4v dpfifo(
	.q({q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.source_valid_s(source_valid_s),
	.state_0(state_0),
	.data({data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.counter_reg_bit_2(\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.counter_reg_bit_1(\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_4(\dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_0(\dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.stall_reg(stall_reg),
	.dout_valid(dout_valid),
	.empty_dff1(empty_dff),
	.source_valid_s_process(source_valid_s_process),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n),
	.out_ready(out_ready));

dffeas dffe_af(
	.clk(clock),
	.d(\dffe_af~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(dffe_af1),
	.prn(vcc));
defparam dffe_af.is_wysiwyg = "true";
defparam dffe_af.power_up = "low";

fiftyfivenm_lcell_comb \dffe_af~0 (
	.dataa(\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.datab(\dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.datac(\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.datad(\dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.cin(gnd),
	.combout(\dffe_af~0_combout ),
	.cout());
defparam \dffe_af~0 .lut_mask = 16'hEFFF;
defparam \dffe_af~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dffe_af~1 (
	.dataa(stall_reg),
	.datab(dout_valid),
	.datac(state_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\dffe_af~1_combout ),
	.cout());
defparam \dffe_af~1 .lut_mask = 16'hFDFD;
defparam \dffe_af~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dffe_af~2 (
	.dataa(dffe_af1),
	.datab(\dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.datac(source_valid_s),
	.datad(out_ready),
	.cin(gnd),
	.combout(\dffe_af~2_combout ),
	.cout());
defparam \dffe_af~2 .lut_mask = 16'h6996;
defparam \dffe_af~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dffe_af~3 (
	.dataa(\dffe_af~0_combout ),
	.datab(\dffe_af~1_combout ),
	.datac(dffe_af1),
	.datad(\dffe_af~2_combout ),
	.cin(gnd),
	.combout(\dffe_af~3_combout ),
	.cout());
defparam \dffe_af~3 .lut_mask = 16'hFDFE;
defparam \dffe_af~3 .sum_lutc_input = "datac";

endmodule

module cic_a_dpfifo_s4v (
	q,
	source_valid_s,
	state_0,
	data,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_1,
	counter_reg_bit_4,
	counter_reg_bit_0,
	stall_reg,
	dout_valid,
	empty_dff1,
	source_valid_s_process,
	GND_port,
	clock,
	reset_n,
	out_ready)/* synthesis synthesis_greybox=1 */;
output 	[22:0] q;
input 	source_valid_s;
input 	state_0;
input 	[22:0] data;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_1;
output 	counter_reg_bit_4;
output 	counter_reg_bit_0;
input 	stall_reg;
input 	dout_valid;
output 	empty_dff1;
input 	source_valid_s_process;
input 	GND_port;
input 	clock;
input 	reset_n;
input 	out_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \low_addressa[0]~q ;
wire \rd_ptr_lsb~q ;
wire \ram_read_address[0]~0_combout ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \low_addressa[0]~0_combout ;
wire \rd_ptr_lsb~0_combout ;
wire \rd_ptr_lsb~1_combout ;
wire \low_addressa[1]~1_combout ;
wire \low_addressa[2]~2_combout ;
wire \low_addressa[3]~3_combout ;
wire \low_addressa[4]~4_combout ;
wire \empty_dff~2_combout ;
wire \usedw_is_0_dff~q ;
wire \_~2_combout ;
wire \_~3_combout ;
wire \_~4_combout ;
wire \full_dff~q ;
wire \valid_wreq~combout ;
wire \usedw_will_be_1~0_combout ;
wire \usedw_will_be_1~1_combout ;
wire \usedw_will_be_1~2_combout ;
wire \usedw_will_be_1~3_combout ;
wire \usedw_is_1_dff~q ;
wire \empty_dff~0_combout ;
wire \empty_dff~1_combout ;


cic_cntr_kka wr_ptr(
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.valid_wreq(\valid_wreq~combout ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_cntr_0l6 usedw_counter(
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_0(counter_reg_bit_0),
	.updown(\valid_wreq~combout ),
	.source_valid_s_process(source_valid_s_process),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_cntr_jka_9 rd_ptr_msb(
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.source_valid_s_process(source_valid_s_process),
	.rd_ptr_lsb(\rd_ptr_lsb~q ),
	.GND_port(GND_port),
	.clock(clock),
	.reset_n(reset_n));

cic_altsyncram_1lg1 FIFOram(
	.q_b({q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data_a({data[22],data[21],data[20],data[19],data[18],data[17],data[16],data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.wren_a(\valid_wreq~combout ),
	.clocken1(source_valid_s_process),
	.address_b({\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.clock0(clock),
	.clock1(clock));

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\low_addressa[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_ptr_lsb~1_combout ),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[0]~0 (
	.dataa(\low_addressa[0]~q ),
	.datab(gnd),
	.datac(source_valid_s_process),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.cout());
defparam \ram_read_address[0]~0 .lut_mask = 16'hA0AF;
defparam \ram_read_address[0]~0 .sum_lutc_input = "datac";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\low_addressa[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[1]~1 (
	.dataa(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datab(\low_addressa[1]~q ),
	.datac(gnd),
	.datad(source_valid_s_process),
	.cin(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.cout());
defparam \ram_read_address[1]~1 .lut_mask = 16'hAACC;
defparam \ram_read_address[1]~1 .sum_lutc_input = "datac";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\low_addressa[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[2]~2 (
	.dataa(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datab(\low_addressa[2]~q ),
	.datac(gnd),
	.datad(source_valid_s_process),
	.cin(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.cout());
defparam \ram_read_address[2]~2 .lut_mask = 16'hAACC;
defparam \ram_read_address[2]~2 .sum_lutc_input = "datac";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\low_addressa[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[3]~3 (
	.dataa(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datab(\low_addressa[3]~q ),
	.datac(gnd),
	.datad(source_valid_s_process),
	.cin(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.cout());
defparam \ram_read_address[3]~3 .lut_mask = 16'hAACC;
defparam \ram_read_address[3]~3 .sum_lutc_input = "datac";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\low_addressa[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

fiftyfivenm_lcell_comb \ram_read_address[4]~4 (
	.dataa(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datab(\low_addressa[4]~q ),
	.datac(gnd),
	.datad(source_valid_s_process),
	.cin(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.cout());
defparam \ram_read_address[4]~4 .lut_mask = 16'hAACC;
defparam \ram_read_address[4]~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[0]~0 (
	.dataa(reset_n),
	.datab(\low_addressa[0]~q ),
	.datac(source_valid_s_process),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\low_addressa[0]~0_combout ),
	.cout());
defparam \low_addressa[0]~0 .lut_mask = 16'hACFF;
defparam \low_addressa[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~0 (
	.dataa(reset_n),
	.datab(gnd),
	.datac(gnd),
	.datad(\rd_ptr_lsb~q ),
	.cin(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.cout());
defparam \rd_ptr_lsb~0 .lut_mask = 16'hAAFF;
defparam \rd_ptr_lsb~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \rd_ptr_lsb~1 (
	.dataa(empty_dff1),
	.datab(out_ready),
	.datac(source_valid_s),
	.datad(reset_n),
	.cin(gnd),
	.combout(\rd_ptr_lsb~1_combout ),
	.cout());
defparam \rd_ptr_lsb~1 .lut_mask = 16'hEFFF;
defparam \rd_ptr_lsb~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[1]~1 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(\low_addressa[1]~q ),
	.datad(source_valid_s_process),
	.cin(gnd),
	.combout(\low_addressa[1]~1_combout ),
	.cout());
defparam \low_addressa[1]~1 .lut_mask = 16'hFAFC;
defparam \low_addressa[1]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[2]~2 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(\low_addressa[2]~q ),
	.datad(source_valid_s_process),
	.cin(gnd),
	.combout(\low_addressa[2]~2_combout ),
	.cout());
defparam \low_addressa[2]~2 .lut_mask = 16'hFAFC;
defparam \low_addressa[2]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[3]~3 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(\low_addressa[3]~q ),
	.datad(source_valid_s_process),
	.cin(gnd),
	.combout(\low_addressa[3]~3_combout ),
	.cout());
defparam \low_addressa[3]~3 .lut_mask = 16'hFAFC;
defparam \low_addressa[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \low_addressa[4]~4 (
	.dataa(reset_n),
	.datab(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(\low_addressa[4]~q ),
	.datad(source_valid_s_process),
	.cin(gnd),
	.combout(\low_addressa[4]~4_combout ),
	.cout());
defparam \low_addressa[4]~4 .lut_mask = 16'hFAFC;
defparam \low_addressa[4]~4 .sum_lutc_input = "datac";

dffeas empty_dff(
	.clk(clock),
	.d(\empty_dff~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(empty_dff1),
	.prn(vcc));
defparam empty_dff.is_wysiwyg = "true";
defparam empty_dff.power_up = "low";

fiftyfivenm_lcell_comb \empty_dff~2 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\empty_dff~2_combout ),
	.cout());
defparam \empty_dff~2 .lut_mask = 16'hEEEE;
defparam \empty_dff~2 .sum_lutc_input = "datac";

dffeas usedw_is_0_dff(
	.clk(clock),
	.d(\empty_dff~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_0_dff~q ),
	.prn(vcc));
defparam usedw_is_0_dff.is_wysiwyg = "true";
defparam usedw_is_0_dff.power_up = "low";

fiftyfivenm_lcell_comb \_~2 (
	.dataa(counter_reg_bit_2),
	.datab(counter_reg_bit_1),
	.datac(counter_reg_bit_3),
	.datad(counter_reg_bit_0),
	.cin(gnd),
	.combout(\_~2_combout ),
	.cout());
defparam \_~2 .lut_mask = 16'hBFFF;
defparam \_~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \_~3 (
	.dataa(\full_dff~q ),
	.datab(counter_reg_bit_4),
	.datac(\_~2_combout ),
	.datad(\valid_wreq~combout ),
	.cin(gnd),
	.combout(\_~3_combout ),
	.cout());
defparam \_~3 .lut_mask = 16'hFEFF;
defparam \_~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \_~4 (
	.dataa(empty_dff1),
	.datab(out_ready),
	.datac(source_valid_s),
	.datad(\_~3_combout ),
	.cin(gnd),
	.combout(\_~4_combout ),
	.cout());
defparam \_~4 .lut_mask = 16'hFFF7;
defparam \_~4 .sum_lutc_input = "datac";

dffeas full_dff(
	.clk(clock),
	.d(\_~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(\full_dff~q ),
	.prn(vcc));
defparam full_dff.is_wysiwyg = "true";
defparam full_dff.power_up = "low";

fiftyfivenm_lcell_comb valid_wreq(
	.dataa(\full_dff~q ),
	.datab(stall_reg),
	.datac(dout_valid),
	.datad(state_0),
	.cin(gnd),
	.combout(\valid_wreq~combout ),
	.cout());
defparam valid_wreq.lut_mask = 16'hEFFF;
defparam valid_wreq.sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~0 (
	.dataa(counter_reg_bit_2),
	.datab(counter_reg_bit_4),
	.datac(counter_reg_bit_3),
	.datad(counter_reg_bit_0),
	.cin(gnd),
	.combout(\usedw_will_be_1~0_combout ),
	.cout());
defparam \usedw_will_be_1~0 .lut_mask = 16'h7FFF;
defparam \usedw_will_be_1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~1 (
	.dataa(\valid_wreq~combout ),
	.datab(source_valid_s_process),
	.datac(counter_reg_bit_1),
	.datad(\usedw_will_be_1~0_combout ),
	.cin(gnd),
	.combout(\usedw_will_be_1~1_combout ),
	.cout());
defparam \usedw_will_be_1~1 .lut_mask = 16'hFFFE;
defparam \usedw_will_be_1~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~2 (
	.dataa(\usedw_is_1_dff~q ),
	.datab(\usedw_is_0_dff~q ),
	.datac(\valid_wreq~combout ),
	.datad(source_valid_s_process),
	.cin(gnd),
	.combout(\usedw_will_be_1~2_combout ),
	.cout());
defparam \usedw_will_be_1~2 .lut_mask = 16'hBFFB;
defparam \usedw_will_be_1~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usedw_will_be_1~3 (
	.dataa(reset_n),
	.datab(\usedw_will_be_1~1_combout ),
	.datac(\usedw_will_be_1~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\usedw_will_be_1~3_combout ),
	.cout());
defparam \usedw_will_be_1~3 .lut_mask = 16'hFEFE;
defparam \usedw_will_be_1~3 .sum_lutc_input = "datac";

dffeas usedw_is_1_dff(
	.clk(clock),
	.d(\usedw_will_be_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usedw_is_1_dff~q ),
	.prn(vcc));
defparam usedw_is_1_dff.is_wysiwyg = "true";
defparam usedw_is_1_dff.power_up = "low";

fiftyfivenm_lcell_comb \empty_dff~0 (
	.dataa(\usedw_is_0_dff~q ),
	.datab(\valid_wreq~combout ),
	.datac(source_valid_s_process),
	.datad(\usedw_is_1_dff~q ),
	.cin(gnd),
	.combout(\empty_dff~0_combout ),
	.cout());
defparam \empty_dff~0 .lut_mask = 16'hBEFF;
defparam \empty_dff~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \empty_dff~1 (
	.dataa(reset_n),
	.datab(\empty_dff~0_combout ),
	.datac(\valid_wreq~combout ),
	.datad(\usedw_will_be_1~3_combout ),
	.cin(gnd),
	.combout(\empty_dff~1_combout ),
	.cout());
defparam \empty_dff~1 .lut_mask = 16'hFEFF;
defparam \empty_dff~1 .sum_lutc_input = "datac";

endmodule

module cic_altsyncram_1lg1 (
	q_b,
	data_a,
	address_a,
	wren_a,
	clocken1,
	address_b,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[22:0] q_b;
input 	[22:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	clocken1;
input 	[4:0] address_b;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

fiftyfivenm_ram_block ram_block1a0(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk1_output_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 23;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 23;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a1(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk1_output_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 23;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 23;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a2(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk1_output_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 23;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 23;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a3(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk1_output_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 23;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 23;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a4(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk1_output_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 23;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 23;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a5(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 23;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 23;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a6(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 23;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 23;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a7(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 23;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 23;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a8(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 23;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 23;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a9(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 23;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 23;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a10(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 23;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 23;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a11(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 23;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 23;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a12(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 23;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 23;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a13(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 23;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 23;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a14(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 23;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 23;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a15(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 23;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 23;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a16(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 23;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 23;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a17(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 23;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 23;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a18(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 23;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 23;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a22(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.clk1_output_clock_enable = "ena1";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 23;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "clock1";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 23;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a19(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 23;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 23;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a20(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 23;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 23;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

fiftyfivenm_ram_block ram_block1a21(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(vcc),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "cic_cic_ii_0:cic_ii_0|alt_cic_core:core|auk_dspip_avalon_streaming_source:output_source_1|scfifo:source_FIFO|scfifo_vs61:auto_generated|a_dpfifo_s4v:dpfifo|altsyncram_1lg1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 23;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 23;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

endmodule

module cic_cntr_0l6 (
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_1,
	counter_reg_bit_4,
	counter_reg_bit_0,
	updown,
	source_valid_s_process,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_1;
output 	counter_reg_bit_4;
output 	counter_reg_bit_0;
input 	updown;
input 	source_valid_s_process;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \_~0_combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;
wire \counter_comb_bita0~combout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h5566;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A6F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5A6F;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(updown),
	.datab(source_valid_s_process),
	.datac(gnd),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h66FF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(updown),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A6F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule

module cic_cntr_jka_9 (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	source_valid_s_process,
	rd_ptr_lsb,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
input 	source_valid_s_process;
input 	rd_ptr_lsb;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(source_valid_s_process),
	.datab(gnd),
	.datac(rd_ptr_lsb),
	.datad(reset_n),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'hAFFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout());
defparam counter_comb_bita3.lut_mask = 16'h5A5A;
defparam counter_comb_bita3.sum_lutc_input = "cin";

endmodule

module cic_cntr_kka (
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	valid_wreq,
	GND_port,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
input 	valid_wreq;
input 	GND_port;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~combout ;
wire \_~0_combout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~combout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~combout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~combout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~combout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~combout ),
	.asdata(GND_port),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(\_~0_combout ),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

fiftyfivenm_lcell_comb counter_comb_bita0(
	.dataa(counter_reg_bit_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\counter_comb_bita0~combout ),
	.cout(\counter_comb_bita0~COUT ));
defparam counter_comb_bita0.lut_mask = 16'h55AA;
defparam counter_comb_bita0.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \_~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(reset_n),
	.datad(valid_wreq),
	.cin(gnd),
	.combout(\_~0_combout ),
	.cout());
defparam \_~0 .lut_mask = 16'h0FFF;
defparam \_~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb counter_comb_bita1(
	.dataa(counter_reg_bit_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita0~COUT ),
	.combout(\counter_comb_bita1~combout ),
	.cout(\counter_comb_bita1~COUT ));
defparam counter_comb_bita1.lut_mask = 16'h5A5F;
defparam counter_comb_bita1.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita2(
	.dataa(counter_reg_bit_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita1~COUT ),
	.combout(\counter_comb_bita2~combout ),
	.cout(\counter_comb_bita2~COUT ));
defparam counter_comb_bita2.lut_mask = 16'h5AAF;
defparam counter_comb_bita2.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita3(
	.dataa(counter_reg_bit_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\counter_comb_bita2~COUT ),
	.combout(\counter_comb_bita3~combout ),
	.cout(\counter_comb_bita3~COUT ));
defparam counter_comb_bita3.lut_mask = 16'h5A5F;
defparam counter_comb_bita3.sum_lutc_input = "cin";

fiftyfivenm_lcell_comb counter_comb_bita4(
	.dataa(counter_reg_bit_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.combout(\counter_comb_bita4~combout ),
	.cout());
defparam counter_comb_bita4.lut_mask = 16'h5A5A;
defparam counter_comb_bita4.sum_lutc_input = "cin";

endmodule
