-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
YdELmdAgs8XCAD4HDn23GOqYs6jRTAgBI3SuRbMWfERlEfJYrVjPuAuSuXMlzuaK
HnZlAnf8guBBlY8J69nyZrxVV5QvJ/sLbPtfrY/R66P0jY8kqeK/BNysIj+mwqKO
wO/Xs5hI+kCKMtQjzrLY6QmM2i65BvzYKh51W3Bdf5U=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 3680)
`protect data_block
VVnWKNiWQ3DBDrkUBMJ0iya2BPUfgi3/8I3tnQu+WfBsfRyqzv2BeiehAxi3DYnw
KQRqm5/Et+9FouCvheK6FM8QXVEufHouddOIKOEzCD5cNvpSF4mRuzWr4iXoSCxA
ZexPmUpk6L2PCbf/LpKZvTpNmaqgWLWEobaF/9ZL8/cA5Q2imPT8p539N8mbH7RJ
j/v9bwjF6iqtd1CqpnCHAH9251n5HzgpMPPK/y9wk0+6hEKufm0BilQuH4hDtKa+
AsYmIp2/HgQ6RZgWI4rRV76tMKXcDkuBOjEUulqtvgEmI+VvHDtmMxGYF84zqp1M
+bU2NfhUEgrDzcoDGoDotEXnY8DUFyLg//hcKWFLBFpv6Qa46ssAZ5Mt/UFxA0Ox
BSuRwj6aY035yCDyheG88nhwmUWyqfomwfVIlWaCh0wcl9gTPyo3R8nKY2EP9MA8
Ma9STtDuCLepdNRebWYFBghDh8qDIzDq3vVMMvvIO/I3RxllqNgogkbSpBPJvtVY
7/b74ZFQjiL2S5zTrKOzWbWka+yoSb0cgcMzn6CaNovWvGrZ27/FLibHHLuEC0Fo
M0ye7KRylVZtpMbEEzZX5t4I3c+rushB/HUBDvrtNqDrJ9KGfLkS19vPMXw+jWNX
8B5+4d1S8SLxZHyO9m5AO51oYGST2HWfZzwtuquczJhmxXPgBUGAgLYRBcYPgIzi
6zAwnLrjQTDFUUq8CssI+xqhJ2mlakUKkaZddYdmOyHW9J6a3axt3yB/NbpE25+o
HkOvBsh1Q7s4myd+Jou1pblFBzmPJi6vm9Jd+eIy5/ITCfBy4O+4Q1O3vqL6xcUR
E+rns1NyQPBZyIXNR4Eu0VHutBN+TWmLcj1uuJR1cv8uTFtWod++UjDhoprptB0V
OjnEOAsbh0b5xmMn5inHuAKc26j/mXwZpVcQL71093lmw7x5I0kO9Fc5t2vr3Epn
yFv3wv/s2PfffZ/TdRw6Pt0AnvmRBKWqmmdEdMExxaLDjlsVStx3qbthnN090b4R
m1RSH1B0yN5t+rLblWI+8oYh+H0Wd7mgqjQPjllP6YgnmZNIfMw/jYbItlX7uzMW
yNJfaN1BGLRDfizrU+hKHrhUFERcgEZjw3OOuKaiCRj5dfW7nVjjCTiuw5KMxsVI
KLtC6af4jeDisjSHlV7H+FgkfXornIlpylR2omNtabEZgunv7R65twKgaag+qjWV
kXaJB3MSZAAlsbGyac+JdD1Jsy55c/IXcewuoP3JZFJMHEmpSQb6KYY0oUIxv4H9
bBMDwccmdDLK+hJpi29ySKJKSmRXhWhmQIyE4+G9ySPRQLlwgYG7olIOay/JQskc
YZWwL7SycjK+5Pu/MPppZ4HcygrpKU+1+t82YFCUKh1WK3LKUI1FpTN0ACAVkl1k
fvUz7cGQ/6vUJDzt86ADL4yIUTv62+9iwrM8AUula4Nql5Ze/taZIQ9gwWYHW+JT
bf8kEa7zqaMuC23BvoU7FFYTOCAtrtOgSnlPWgqGJLh9RYAELXCKZcdqBwUg0ts8
Mp7aKca1mkTasf7SHjWDIXdo5ZuD582GUBQ8Xvnrccu3t7asTzm0F8Z/yxLHGAd+
OixR0hPOtC0uRhsnKhekqM3QjIl/oqGSX4GvvsI8K+7Als8ZeyQVIUO8RAS1Y3lR
QMcJF4CI1PweYT5AaGj1aj1e8puxkQYEIYySKBugoFnGf8QsjyjEXkH9B+HWOvCh
FUiPZhS1VmM6Zhv6icq11a571ScsnEyXwYPKKsAhgOyH8oLjFAh4JuWj+wDJRASj
An/T1udhxvSmZ1J0NJ9Jirm5sfdlw+wTje6namjlGOq6DpoPfqziNJtrfthStM/u
ZmKP+zFkHG1WyrSPGvBVSqMKnQpehO8BJMd0RhiT2yjr0ChXTzQTp9IoYFJC6vZD
qrtg/ZJAQq5rk9DN4qHnEHrHmwNTE2AtYt6y4Ts6KBSt7+8jVntPnGQ81AIKymeC
Ye40jr8+F+At6sJAcmnvNVnr1F9DGO6GdjDsd4WgTsJy4zWcrAbjNVyJ3/tL+X4z
msKVaQYRAy1Nhxlbc23afzO7Ou/k9ZieFoJrlGmzIZb1FFMDZF18ZbVRGZPMNAUU
/UHJ87rE/LABG5qz3BohCUL8ApnbE0K3zZYTxpprACY2FPCnAgBOCOqUoF5CqmrL
uUroHR+2vB22/EPjsHdw4eHtYGokxKO0SDoNJopgwNSsWFegNPj/kte8WLghSV4h
gQ9cfnZIjjuxtlDH6+blA6E2XBUhi1PxdB1XQhe8JBMxu3ybXK+RpK3dDECV7E8D
IaJDjo3F6XxNVFyOrB6lbs7X40JGrv9d/0pzqSZ9N63+eCyGPYqAvTRgELtZDSGM
Rj2pN1mjHGkIzGxQLiM2+Ol/Mb7OHMwNV7OSiMHJDgLaKA/E6ONEqREUfCkWWhV3
Ed1HgJPjEImYxUlBU0z7KGoM/QV2xHATDApq4KsOT/pTZHWDkjqnhHGx6xYE9xkM
XMsdUPMKKdV/ywq1Pcmq1TK6n86ROzEUMzwTUNlWSyX9HIFM3sYXQ9r1WRfpzoXc
ElD93J6gxV5pQErEXBMchFgbwkvYPzz2TzV3b7G8xf3hkgYtl5iX7s1BfoCtpgls
y0TJoG6Py4eD9mai69qm3WpH+cJUALcH1niSuf/QCObojA+xwRnAZOsaxx6YXbee
wUaXTgEgfrGNo7/SRFe+tSH83EVypFzpKaUqDggrHQ2e85Tsdhi15QNVVb8NRIlI
K/Uc8L7QXpWQLuhF1wVLck7ZrGJL7j62cf8Wu7hegSn66AjHeUeeRUfaLRkIOJPw
BE/gMetzc9pcuLx/Xy5UuVWuvKVH0ToJuoY8n0y2yZN6Fa+oUkUTFWx3guJb6MeN
qTXZo/LqZEVPw/x2wKZdt8zuiy9Bq1qzHduiK0D3Y800TgQ2WNps5ULiwCYkjWkJ
Hsl3nl2knOdH+mq+DVpS/V+SY8J2mu0+0GG97fzjvOA/Zd3JJ1rIYIYRSRtM2R8W
FPk5apxevFSnJ9+nQdr+mSGDRvOl/sxW4BvbQJcTsWoAVDsmCQ5pVh7Jfi05swti
OMmbi9wgFb7RBxsyenYzWX9LT+scGU3fFctABbmeMKbWp7EB3uAH8LQyojp+1w6t
QCF5LZd+LD2CcGhIpOAU9XHXi6psUJvsnrSmuTOXKL2Y7gZcR5PohTxeYhEYeLgb
TRGdHpcfYyHonciUupnahei7d/Io1zTEmSRfzZsUuvUqnPoG/jZIt1Etg+rktY+5
pG2fwa7613xppLP3tGilZLQoChfqN57VwUyQpVyqRwh88q8/GHUD4fWUhjYKssiz
FhLkte1o9CLi3QjHcaMH4OzbXlrfilP4JzCJmAWkMzoATRv+92caP4ITVp/HeF5p
81QU1IVZvOFI24A/mCpHvAGCWATYNoXf/EoFVa4COXZf+CXgxenEdYXxePh1jEYc
4ysU9PT+N146Xzn/eShMgu2ScRxE6mJzAqS22Dz0ROlGCEED9gO3KR2JUgNgb3zt
u/p1xgYeJm+DrGHKwkNJZ++Mirdq414JD+T9714nMkkSDWxK+3Ama+avovx+WjjV
9V7InOXRN8W8yTj/g5LohqRoe2fY+ws7KAmGMCDZkKMOFemTKUDvbLvOEgDhVHYy
rT2iYa6qmUSNyulgEO18TB9FREKKcVxSjGBPG14rwTQn91ZFrjLMeruWE0JsktY7
H5yNNg9LYl0wsyEqQGm6Pbafuj0MOUCi+oRWmzg75ozrgPQEeJ8VcCH7e1iDyGmE
WNoKrOqyj28/rhV0xHQFwkN+zWq169QgJbdsZWmCGljsvXSZx2Wm1uyueZsq1Ix2
Lml2wvL+fNqB8d8YXR/KGiqvjixJolPzJcyFT/EPqlZqpU8Y1T1t50MoTpdAWKxQ
uwlSIGf67AOuX3PLw7mGKuXY2HEuhfJ6qEzBfgvvgNY6kL00aMmgp508vMEhiEdz
b++MsZTNs68UskgvO5VFXYYnvOxF7v/RuJ1/1LbeXgHY1EeNQOAzJ+vlDdsU3w3b
mCRZgIzS8cSOL7VsRrJ5BKn5zQ8m01oq2jIxjkIvhsz64/UUbX4cpWAmZa3TX9HQ
AvTkSn160z23UjZ/vKGWF87JupdVw8EE0wAuRNnDQIT561iZWNCIJpCHxrVeo+3T
llW5vGnAwXtl1c+qia6iffHiuWPRklvsp9jLlvxyhWIIswv8NDSx/Lefn21XEMRY
9YrJ1C4xHv+p9ZpVKpHxerE/Dz2yyNaOu5pXvA1tkCtANGhJQXGMOkbWkseJRLob
6iIGQyzB9NeIflzgcGEH99Lz9uHdN3s27evM/0lprBtIYuXs4tRK9b7sZymxil+c
k3lO+E5tNoP7Jf5AaFJqmKmAUDRz6OOl6IZhcAmGDquoQh+bl4XVQclUL/4h0fIX
dI/e4kqraMZ29pv3qZAszxxXuS0mQ1S5W3ffiVS1Et66VU4FmuWYNgoQTvwBp6hy
0z+hxyijGQe78tD+Kmndrqa2ZrOqjX4L7I0DLbmM1hUYsH6SQL7p4N0cdeAmMAgn
BxXFU9RInLxF4Uhq0PYiS5NzFte+J/Lp0MrlsJwNnTisS3tmhcw2u1LmJ2sjNzGY
XHo8/QTgcNDpobwTuH3WLXvBs4f4NBF+KjqF2xXZAdKj0/F1x4DnjkSY9L++UExJ
p0EMjV8ncKR1I7xsPcdEwziBLonSvdBGzbJoXVhu/exaOR8hLjwQSj2TTUrVk2sr
ph8Ma4C/zhM4+N0wZqfigG5WQ8IF+YyfIASzdnpZILgDR5cvIqf6BctW/Tg0LtjA
RIXwbyh0ALjNCF5MRnhQdeN0oX2VR1RIWz9hxUVAs8WyYizmkDICgcliVbbpA1Q3
Is64Dv9qRnhs+2Gmxq+D3dQFTbX8t5/ETb7R9YzRLwM=
`protect end_protected
