// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H8Q"0&ERPHLW,U>=X2E%J$#V-A<SG4ODG(UA;X!"M4%0P0"EUL)5X9@  
HKD5JKB8P-]'V2/C]O%^5LXUQQVD?#.4I57*U'R2OOR0#;;?/V6XRKP  
H4W7I!AEY38"IG\C1=;5.M=Z&K[V@AZGVG#*U/=AC8ME]I6M_[!A*%0  
H8$;Y;WC.VY9 =.N^K E,IQUB9"*R>#Y/G1P$?-_UIJ!M*!S.'(IEP0  
HEWN7(<E+E?@BGYR/2A(TAVL$B?@TL+WSN%S(2LE/%KK$=),*/U!$WP  
`pragma protect encoding=(enctype="uuencode",bytes=20480       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@.B*+K5&HI(K_"F%T90+X +S,LGX0=]A;RN'[4=!2V"L 
@QM"N>NWG?3/V27CSJC,Z8FH.1:+B3$AW=<BS2WV^&<, 
@MT$*E![J4L+M_M !$DY8.WIROH"L#4MPN@'31XOWX%( 
@<3XUFXVU,[+J<JY"5W9?'6^5SVNGTH&72 'UI419%Y\ 
@<!/9Y&"%O[!PJFU.?!W-L5_Z@A G\R0=8@6=E-DJR(D 
@4N3RN6NAX,G@JCP1V:V041_RYDI;KTIEO1"* GOSBT  
@S*>O@< 9.!5!2N[] RC1+O(G?IL.#C9I/\6QIQ)4HVX 
@0C%%/5H?CS*8RPX\(RGQK2)7I"M!!VEZO'[L.@V*5%, 
@F!2=B02!_]QK:FH3>S2)-%._IRD!T<8C!9LW")+_*!\ 
@L<=. KXHR>X8PCP3DQYXKT;[Q(13+EYG!2(G@6/%Y9< 
@'\/IS[K_>U%%TM-&P* H? -X27F'(1#'PD(JCW?DDS@ 
@8=FJVV-8;\SFC0X>B2 B< ]HN=<V8]OV%+WP@.*@L$\ 
@2LPH/VA>>&B/K\[,S?ZH!R*ZVPDAV.4Z2OLV$CK_4M$ 
@E#J[83FU'5-8_U_86>?@AZJ4)]^!A=D%Y%NL=I(!"7T 
@T[XD14L3V.?JRY$E#:>".IRM@IC,*J-6J66",)>ZDRD 
@^862/D:FD:[IE]0'5#Z':J;&\ 0':C+8/61*+OG,%MD 
@8JO@N+-Y%D,3POT[N(D=MKU/FN>&4L-#++:N\UD(FKP 
@[C;'.W^WH@HOF"IE._,::C[+!]HJ*L_O(A(X<7C'!P, 
@S+V*?T3YSV"L>] ZE-?844EO6_:%08AY6#I9OI W$ P 
@#B+=9*7&PK+9<-<IUCEK!L.<MLGND')U!SUQSVEBT8, 
@>PG.Z^"9*]&4MQ ?M;X&(E1)Y*7JPI PI14[< ]T&%( 
@N8AW>$F>!:ZNSEU)DGNA0?SNTU[WVU@M@<,0$@'VN8@ 
@UU"SP2XJ1T.0 N'&$[@PFC_0Z>S[7PHEDC?1UI@9X78 
@G+@>0G-709:9]:XR"M?.@C0DGL8G<H$P-=-<7;"?!T< 
@L?;T*<%<A2Z[7P)<[4,H4_LQ\S*0K1S0;'8@Z!!> 7X 
@9&2:C'VAMOF$3%C;D5_XZ=6W@0%Z%NMN.8ZO-&QZSJH 
@0![NL@]I3+&DO#]:_E'?PS31Q<WD0D3351/GTDKO6"P 
@4U2;3>?UO';]RR7XMK-Q4A4:G]J=\:H=[Y)SYSH 5I$ 
@R@RAW$H*,#C"A6>\PB<4QA11* MX8^*[*F\8!G^(](H 
@\<5N&AM6+0VER>Q:!(? T^4;GC6FJ6#7Y3 ?P.)POAL 
@X;F':AA6V+B7%/R))?^VG7IC\2ME:0K:@ =$3#.>AV\ 
@AT]J,[?-IF1K ;&#/B+RJ$<K_^C>&K0:[K"(_]($E.  
@))HHHJ=#\(O2OT7JS.1I7P.69<=:0\%N*I0.N,8I!VP 
@G>? E*7 )^#W9<T8AMO(<U@_<<4I,1IV!\^K7>CAY[0 
@$^6V#_GGLH5AR&:L5V+WTQ-@&N#]^9+K; %"T]3+:G  
@31C_9V&O3PS +Z,[MIT+79[Z0P7/)!*-@>BL2PS!G/< 
@74XZ(J[3OL&X=J?]]9T+5(TX" M2* /; H?W>G[;X"0 
@&2K4\.OJ[:7CR&[5_<ZPW)XS\TVU79G\QB_X7S"<-PT 
@F=;1'H!1W7VEG/F6&>6/EO4E88[QX+N/W#!1:ONVS1( 
@/90FP VRS3LZ#I<(&U6^9SWBM$:C<#7<"9;",TTM[:0 
@-FTCEDVZ:!,_)-$6EYNI'Z:O4$G1L].A==(.RZ?SQXL 
@3+U1-<6^/%3"R8.6_11C]'P&RN*ER$#Y&G]P,2.W6+P 
@I!>-<G:<ZPNW.G,+-'-PZ >_<;A$REK/?GU_G.!L]_@ 
@(SS"_%Z,88C7]6>D6!P& =R-^G@FF80Y4+4#\QF+#@0 
@\"7B>1<Z^[@)!RK0JY9:H\'DN6EIZ/#?MD<4_>6;'_T 
@D6O4]+JUNLG@89)#Z/S5U%@"2A^:E?6L]:U8>^M\FI, 
@HK:$1^G!CYL22]G(,G%PP;PTUN0)_RI9LVPILLY.L7L 
@9(0&Q57S(:0SB1-E899=*B07AD<2W-W_XWAW1;"50^@ 
@@E 3>H/VC_*5V8ZW#"2EOK3'@ATDHVN97L7D>%*SDY  
@1W$S)AJ<*>SP^IVJX:D8VY4TSJ?F*1DL'0; W/A#!.4 
@=7H]\\4J?#.!XA>GR)>8XTS.[-Z8S+H9R;0*Q7RB.X( 
@$AP@X7F'C14:,\(43('<U:6SH[+_3JCGCE8=)+<]M3$ 
@EJ%8.<>ZY5=\^ZHL, 8B!;V0\2\9LJ;AR"!P&WD!/L\ 
@-494/)VY%@/SI1I/;T))W)=&9\?V]9CBO;_)-A[$FWT 
@E+C1[X66TNA]T"D0F7L87'EXG L0>E[0R/98 '7Q[=\ 
@J5+ ;U[W*:=W?PP#-\/[84WB(A.*0X1MJWMPR[YDZ7P 
@:)<Z.NAM:SC MCO6N*LDN/]=<K 26I9,5%U6\^IVXL@ 
@A$0]6/(R*.%8('X/]+-HH/QH6[\$N3-P9A/RD1UW#J< 
@3F7-P\+=Y"EW4I4D<<>MDP8PQNST7MYL9]S5[4J?4S8 
@I;B%JLPT6S] TZTW:1"4W$(N!Z3X0--R3)1'0>_ ?9T 
@2=SN:,]-/R43'RY^T$,6!SN2*.',*/S!9D\'_+^GM3P 
@!Z57F$(M8NG4#*":JREB@;R@UZC>Z*#([Z7>:BB9^_< 
@:QS5@ \AJHC(P=^/I6HJ+1%3Q),I#S!%H(EFSGHB*G0 
@<? ?]L OMF';/P4,/9?_[]NI'F3][^0XA? #&R2#K!@ 
@:0S4TP+A]T<U3NZQAL=%L;3DRCN1691/>T,53,8'C=\ 
@.40V[.T-26-,*@$<D9N^:)5(4ZG9TMO$.9SQS<K:=8T 
@<I\SCM2?<B?'&Q*U! %AF/4C*C'/8I@40/M*82\Z[C( 
@Y5T/#<;<9ULV/SYR63$0PA[Q-O"-$[SDWN>1YQ97SNP 
@ZAB.U-;[\IQ9:?;H.^^7;/\MAK]FTI],$QLY!P,?PAP 
@(ZYI8W8PR[T'7Q3]F89-T:/ ?@%BE$=\M?%B8NE%U%\ 
@(\$,]1'X?5YT1A*C2EP.?<M[\X=_^^) @+U2O!$'[^$ 
@<,"OGP(_U*$DJS0X0!U#+C1_/ (VDW.!YI:':4E0-:$ 
@.G"QYAI$W(G^(\]S=Q1'ZR8=[I-S??K1 4G?G+H8%+\ 
@\M)ZQ.'YJ,W7?;+CR8/33C]$,$!N>F]6!A4)1M 8FFD 
@E+1)Q>9=JH2_#BY!63OJSY'?R>TRQ5K!B38/B)!IX.$ 
@>]=LU:29M!IM:4_."[XCG%.SXK*^SUU]Z+U>E[KELKL 
@+B\]K(AI D]?4*O@BVIMFN:B]5!U28;_RS%;^\L6SQ8 
@SK:6*SJDB>M@$N8A".E_SOIT3 %-@,."!/-;\_@M(Y, 
@6S2>L_L?6$6:X \=HW#\G4-=$2!CBS]C!.BP*4$^L-X 
@Y/BGPE]O<S!PS$2!?GV$[/]?,IG 6+'-'L7C.I#O]3X 
@2"]/T]-[:J.5H <5!**392R<D=7TVLKF:U:TK-^+QBH 
@HA,[&P+U9DQ?TK[@]O3RN>JF=VXHH^53]'J^L6?'&[4 
@ ^QD_$>ZOJIF?,<98PC!C<W?JO833\S5]T#BT;)>4G( 
@V'+FRL>N!"V![J@+ZT#$AX[J8_L]!H-G ,[W@Z9KWWT 
@+"WAHP7+U:UM8RB,]4H+\/I4GG?HXT?6P8[K=@/+7@P 
@0O8'Z\L$HK+#UZF/#LBUSR+7X.;]PB$=UIOT8?(X[=, 
@]4';5H22,X'2WLSZ,Q&,L+.]7^KA(JM5FEU:3/;\-D4 
@P[_('9A+LPRV:J]4?;+8@.)=IL97V3=<!D<_V@85&NL 
@J?)]><2.?I*74A0UNR M 5R32+QO+_@=L'3TGR"4FH< 
@+.>SX:X0".3R&3A"A?[9O3 W'=LXB_?&L%.> 4_X-R  
@?GX;@E+.T%5XU7V5&J4]%C$E=^<@2]^M,#VU3_4\]D4 
@00K_]*4X-]7<;K&Q:# (RP.>77D(U"AU4AY@OFY:S,H 
@J;"6U--_/,IYJ1%M$6:"N:I(W'P0AK3&(U_.#R&]KL\ 
@S0,?4K0C];L#S&\O;,7Q7W?JH2^#!WIB#O+*"&[W4%$ 
@WX%05.W<F2T=O5"M&[%WJOH<F"V(U\Q&'R -G\5G9J, 
@?\N56UORLC[L5Z["5^#RB$&1]/Z\G0"PQ@KW1DCLY 8 
@ FIB6J\@?GE7,[XHD;]@]V!R%%80Q+%J+SU]V#3.)KT 
@WOXRGV=4P7Q'&Z<<EK?I.P>]C14%ZX)?<'\D5I38$J0 
@DT07%XM\BN!WACRH9,A(SKZH_2N '6$=#")YMS4(NN, 
@3=16WF6\0O),(.^8Q8A:F3H(L@Q!;)4"*$=+8>U*P:X 
@$',8E9!1RA>"KBV>8B]4J,=B7!C7RSOM_V\R-;^:+)L 
@6Z0IJH1-./W 3R\2,M_6@=BJ?5<Z#67T^N*4DH]9PU4 
@68VD=C9<MZ^;:<D *\#;"/J[.0XR?Z_+*02;NG?[%\, 
@W-X&$HANK'/%T'G_Q\KDX@6S/K.OL(6WQ!2TD0;I8&4 
@=(U--(M)/[>GLDU)'1S("0HH'[:SSI"H_%C'%!(#:=D 
@)C *N T158_YM/5>7AWR1ZB$:I$B,;+N:^&>03RT1#@ 
@):38"3L-+52)J%W<VR,'+Z+1^C]^0QA3'E$PLS(5L@@ 
@K'E0TDVNXJ>+<([=8J]"2XHW[F=(W=GN(+//8Y6@#2@ 
@5%,3T*M4)['//3; ;E!=U\P+< /LHP]8>?R\=6^Y?"@ 
@GIV)>HVRFU[]^9KIP83(%A6!-_2METO\PB?A"MY.SI  
@M*312)\X7NQE0YY89NX@"P?BN-\_.B$SB-M 8'!8O.4 
@%*A:^@EAR&%YO]U,ON+.R9;CV7@%_GM<4U9R\F,MYZ@ 
@?D/;9!B/'W+))5]L U(4Z0<44LB0-6N+X%.>GO!KWML 
@/V/' '!86+PN&[$A--,AFCC^!K*22!U0*]/FT3[KGW8 
@%;7MAS [LN3X8D-)G*M)%UU"A<&;?@P =:TJX_CZS=  
@W;C_AUX!-.? BWN 8:@YI.(PMJE*JBKCWBJLD\U#YM( 
@Z\V\O]V"XV1\-Q$.%&Z0ZY2<0J_(\+ZZ1,I3]A&EO], 
@C0%!"'C+&USI97@V(4<G;'\+J7"_$L[2K]Y#P&M- .0 
@MT;]-,,+R&Z<LUM3Q+MJPT($9M>9]-G_$J1P>T E//L 
@[S HI"3V^68A^WFQXW+P!7RBJM6EK[F5Q31_(CRY0>  
@U/" O?JGP#.-"GE$W3)JCQ'G"N=8W4 0/;_7JPSK!A\ 
@C!'H:.H'5&CL_=P03R_C/&+Q"C=/C8@-B+KWK]%PVJ  
@\G >T"T"R(]/MSF@HKC!+W<HW"RO?!KP S<S(^X[<,T 
@A'9,,H,MKX0HZ?$2'MJ & F3B^5NH\4:BMH0]:#( G( 
@D4&[QQ*X<HP/(TG1&?@2WQTA0M*O?>&RC$.DYO9RZ=T 
@,C5^RG%B9WWFYQ@STAG)@$H$\F$.P9X\1'3L9X5"2TX 
@4UY_?S(4ZL]$!QZZ?Y*#NDT:"T:49F2%R(:\XA-_S+  
@CRH@<]1,6':@9UO\7'^J(T'T=W,. ?#;\U%M7%@U/)X 
@;AO8K8W3)_((6J@5X"@<O&L)Y,GXC7M+E]".9LA&%'< 
@"*";./BPQBXH1YB7ZJ;$8I*0"*+ KSF9'MH&Z^Y7EZ$ 
@7E(:03+AXV!<ECA9O8J7Q#;Y]A[G53K(.88-R$"2IX$ 
@=_Y/76!MO,D@A=Y>#K"@Z]3:2P>T%7A(+F3^S0OZP.( 
@OM@V4Z0RFJ5COQIK_UNFCOXM!?*01$6J-@H'J#G:IPH 
@*0MW1;B3=OT$-]/SVMRF[ODELO'Z]N*XL2&]S%NK5ID 
@=--V\/IM;"RJBTQS .0/9U156_W$@F5.-\Z%U3_N,SX 
@0ZJ-IT J5,6/16G/:%=U^9DS<33J(BXOD]P&IJO]ND\ 
@]$4/-& J&A$_N!?9'1"KVEP;,1O!)0>3%T-;XP.#+B0 
@,JPY=.(>K@S!HLK7!M%!^A([]B&8A-L^V&Q& S2R%,< 
@'[-P*\+^ 6C0>9 0G<^@O<LVYKAA%(Z,$F$,6<NK^I8 
@9#-/W5A>9*ZA&X.<[XOXIV85UW5#3F4BL'&"X]5K9&\ 
@QPT6<*"M<1HK>^MP50XGPJWXU#+_=8>+^7($3ACF+ L 
@H00-4/\F?54N1(P]!F?&AY#+-F;.$@PLFOY,[X[^D_, 
@CHE%G'LR?D0YQ=(%]&!7N&;P></CX?U7#6.@\^6&I,4 
@7E;$4SDI%'J-[.'@_2+MTU<$&#O!(W889"$_1%%A>7X 
@F.D*,S1T4V4,3(AU+;%TWFN&J5; PXQ3QX/8&01](LX 
@]U2S:3G#=&3WOK08?\Y0$0QSO2P5U^1%!CIC\Q<M'@, 
@P;- _OU"]=.]MPWZ*<H5U>2HZ\E?0 8;+O18@2.=*X\ 
@N@CP3HA%)]HZDJ>*%%\RT4_0FVS/U7)A5,D^'VR;&]L 
@U<3O.,BI:BF8K@0:PD@Z@U!&T4<HF$K5KN<[$F.B/I4 
@@_2"M5ENKRXVVS%%3LCXD0>S+2%3F(#*YN K)Z/&9"( 
@20S:7O)):\5AYBDA@RB9>R3&5TC"]UJ-B\3,L(OKO-0 
@Z<;*:G)?Z=KXVE9?J$0[&\.Y^ABH50FAW,OZ!QTW\@H 
@3VJPBT ?<W43J_CI*JR@+1S2O1TO=4S"_#T\&:C#*3X 
@%/2C,3FK/TI.N"E3"<B]/G2/3_&S*TP3\4M;HZQ0L\8 
@B321AI4T)0!(^9'2DB)?$3^R<* 9571 C8+*W[O-:FH 
@;;1U6MT>M3:^+:AYM,?$P[,O?Q+R-IYYK'-&+C9(%&4 
@+U3GI8[-0%76I[8+2H3DMP$F7J*=S:H[W.KN&+,TL,( 
@WNW4_87:9/O;.(6W]0"F&&U^*O"B$PG'A&U>^)QA628 
@X)MX?)L9GC4*+QZ3OX/Y?]^;4Z"D^^Z71WL\DD;9 >< 
@"DSG3/6^M;PI.V6MM5<"E)M6K,!'N@022]O-SYQ*P%( 
@7'0GTS'\QZBPD08Y'=1+,A>ER PV?W]VA4*Q1(BQ+D< 
@9M"FS"K7"AYP*MA[OYNZ7JF]+$].WOOU.#"B\ZK$ JT 
@NK8'A\WA;JK9U0>G+/4S]Q.-.(C^(!S8I3)OV7VC.DT 
@[S,RJ2R,S2X>_@!=*L:;SM@_B!]S02*>17;%2Q?7TJL 
@&:E/%7AMWVP>*9/EEG@F*Q@IKIP1\9]$"9V!YA*Q>C\ 
@M;])3KWON-O*;';@V$O6D@R^,T>^@$.^Z +]L&3KZ<$ 
@&5ZVR([;JHWC"1#LQ5/NT$1HOR92CAF %X^=2HHG_)0 
@M&>=Q5+3! N\C4IQL1U"::F<<3<H"]8FI)E$_LWRPM< 
@RH9)4](_'<G,AH,?7^%$MUY:8M/"ZJE33G#2FTM>+@8 
@6!3U/:(^OY<#&C5^>7:SD=&J>-INPSJ_MN2CR&TL)R< 
@2)$'J/F,*ZO3Y_/J9Y\UQ"K<N]\IA.$=6;=H5')CX%< 
@<RD+Y#;Q_)1 ,^N8=<:YLP+59D2-S:-JV+'3;[\>>N  
@=45 ,)KUR3SRAU>F6DH5GFW!E2G4]'=I"L_Z9(P>17( 
@UV.PBKXDZ,A=>/6V"D'\]%D0' L,+RY1(A>CA/<B):$ 
@ ![*V6/9C6KLE:CR<P3UM*(810EYG\[%-Z 5:Q[%Q%( 
@/[%J#_ATO_HTHEH\N5#_^=BX2O_79U6QW6NYJ$](D0P 
@,:,I;B'QY&8!DEK=,B#%%L\DM>/?*\2FC:6:2,60VQ4 
@-N]F[!7"HHW@Q63U9H77;!(..YTK"\XK, 8>KV.%=L( 
@Z*E3_9F6%)V?H:$C=\%D$R+"&GC/3)60B/-$&AN")"T 
@S AM"?**DV?F]P80$KVO+'>]2R00 GGN@!2B[@$HX6H 
@C[.G=AV?;FJ#K]TK0?*I8DI;=0%>'I7L?LXD)Q$&E&0 
@YY&;4%YLT.?_U\L.1WT.HSCH<KF<;:9#+]B7?N0\"E0 
@7H>%E]"&:4:4BM8['1#[4K&J0I#'].@)FX$?ZF19G<0 
@+R 2+HNB^!%WCK 1KW7)8(T=  LGOUH*,GL%<53@0'T 
@5#(W-88^0G#9PDIX%R VX!V67=^CY,L:2(O]*&&A3-< 
@[8N_<97*^BP*'7[\0)RH;J5'R5K^Y"Z![WT59C3@654 
@!;CU#23?-0J$R+TU-=6V_."6?D!*59M[D/;;*HX1,S< 
@2T8\ $^'SY**_XE,81Q80%0[%?O/B^>07O6&&C[4VA, 
@&DZOGS8>[+6R 1/"'JK8(:,-VOK/)T_P[+J@ERI]Z9$ 
@C^7-+<2,"A^F[\C3#!1\CF3&[OE$CXJ0L\IS[/,5WW< 
@TTG.EV7<]JQ4/(!Y1Q+-=T</!*EZ)55E+818#UGN8Q\ 
@]"E@#7C$?W=HTP2B&[V\=5=F]0V'GT:4%Y^PGG'VB!H 
@EJM^8J!^3DD.^%R$=66$0TD<9.*BPU-2=Y99?C*8.[D 
@@NZ*DGU4[,/#T7?'<VE/K/=;PK";4U&(/.BK+J(PBH4 
@+(GP@C?$]_)C.U^2 [5Z^N:*R9J#6UR,Z\&;:*$@VRH 
@FDFA:%SD"!:_46PZC-L5E#A?<L5/L$*H!W10Q1F("=( 
@SY#LH[C[LEU**MN'KY$HGH2>AS'E[K(F#2GV=T4;L[$ 
@&_Z%>7W@;)5("<N>(E2Z6&G[^FLCFOQ57#N*G*FLZHP 
@6W;VQ6K'<"3)5G2NB[8?_ \:?R+&4Y)!N#-T[A[;L.L 
@*E0= 3ACQ4.<N_M\Z2W[A&T<G5 2+<YU&Z./1-5JJB< 
@BMQH<[6Q%RU_^&8,,;UF9YL*T*-%5P+?R%=W9QQ$T0H 
@3T0*AO[&,*,+^2)J3F4^J#VL;);W4A']GK>;PMQG@2( 
@RJA/XC?N<]X3+ZACB@?"?EL;T &-7&-4;?F!&F*J&K4 
@J#0 P2>%(,#\Q@Z*8\W6WTB8,/ ?\4O>D6NKTEW=0@0 
@.T6(+GSO/6\]U>[8N5>N'CP)SO\N""(3]>;;$<@,<>  
@RV0=P1/D8RWG!M&$RPA'^U93&3]VF>8@]E0%3:091A4 
@YF]$-RUXS(@\+[>4((R.*!9 /SM1[0W;2"K3[5]&NP  
@-M$8*&=''^^#E>"9#T45*5U]J=V_$#Q#(@RD]>#4OOL 
@<$THXH=0^0,XR-')WF"O@C)]JWQUQ>3N#+(>6X(Q.LH 
@W''A0'\O%8MCB&#K@S;5;HRI:4!FW( >.4+KSJ(68R( 
@7;5[)H@N5AK4*MZ_$Y&*(=)E4H*53%[R<NOH8.()7ZT 
@<4LXU9+.//ZL17%U#H^*M$ ^?(B=*XMRNL7=-EUT8]D 
@*>=_>9N*PZK6&5@:T%[-MPN9.8[;9%G Q+E7L[D7VA\ 
@YY;.HP'*Q5)I"MW?V\M<:@FCX"(\'PZFQQ@/;4Q^;J( 
@U1_=-2P*B\P]R[@NFX/0Y$=9Q+N\3\*FZ_G8Y YN?:@ 
@;AU79V][Y=M"LV-F0=2'8,KK#+.M*L#8 C&#507^U7@ 
@2<YBZ(6U-XY3)!CQCX"=],IH1A-(:^,P!]@&4MU2:^\ 
@C!4I48==7''3&Y3;#/!(/&EX_EI%;MFL/_K!GLJK\98 
@U_=+[9NC[*T#JE^TD#/V:Y1!+Y_SX9$7)+4 C$#9@V  
@U.@#7LO6K*';4)KN("QAXK'W1(#.P02"ZM^43.Q[E;T 
@ITJLSA"_5Q$ZP=QA [B@'%S2=I$K0A>4(YR&\:/&V'\ 
@8A_I56K&GOKDT?](PDA2&E8-9N;E@-T??E0\2=(Q7P8 
@">X^C\R?C!HSL006UG:"=I]2\J<^7%4)M@-8E!)/9%4 
@K0^SVZ?0!L/QC@>EW1*'="-TO39;VQ/R=8/4DR+^Y.D 
@2IU3/LY6#/#>.<K3.R>,-Y$PTT/7>3QS"+786S6B> P 
@"SN^:C<0A99X[<*L6C]C%*'' A$ZWP130'*47OOIXSH 
@/.G0=<+?3R *N%8[[V?,S979)_O6_+P7P[UIC^DS92@ 
@ZA!+X*9QR"%!XIRUNO1!D?+0%!7]%M<1N=A2IU_21?@ 
@BP0 M\-U=3'(P.,VJ(C@7+\A5-U8N4*9_[2G#)LU%P( 
@G[[%\!]S_9-,IFKPZ01L2F2N$H!4.#EFKRHERJ['20L 
@60Q$\<<6SL=@%7S\U:*TYJ9*.)]H:6<PY$.T,MZRZ>P 
@G8.%V(;.Q]XYF*4B*-O9Q==YY%9>4(>IT2GI>K@>,C( 
@21++4F^_NB,R& PV2$H@M=_IW>.J4]AZ$.@%ORYYWH\ 
@5<8S<64P LD%J3QW!4?K7'Y!RQR[O1,M()MAX\P>EVD 
@7MV/V+/.I]!84,C?\_>NVWOMR%GEU_%!^QX$=L Y@F4 
@!)Q._JAU@V!W2:UI*Q9 D+GLH92L$K.3VZ-KWO.@?ZX 
@RQ?W_[&1AYHW <RF_CLA@^3"-2W@0"__+D@IGF]DW(, 
@IIV+CL<WKMQ]"4(#S<$.D([AVX!)QVM*Y:K62J/[[DL 
@BN'TP+J:_O096+7,WDW<U6P&R.M$/6.1",$)/**YV]  
@-S(A]4[]ZI61>1]\<A:'C(9.&R ,G:IZN9Y^'?_ <D  
@D&OJ>(<C?31I=A1F.4ZCW!ZNF?M\]/MB$*5"+VI+86H 
@B9G3[Y3_BJW,O:??R[+J2AMV$@[9 +C@OZ[M*L\:\ZD 
@9)S3M.H* JZQN]7'P"+2 I;;SG*!Z&=^PX)28CI^SVD 
@M^.O+WT=$C06C108"P):!L\&IJ,]&*\KW#C>LY$!!J$ 
@*WUWTA2D K>>!+LT&;0TEI7IX"MBNH]@X!%#SZN^P<0 
@0VG%\JZVG:N!M!5!+*Z; MD#XT..[/*?MO>[W[ASYH( 
@-PE)J_E/ H U'IG*.H<S]])1),D$J9UIAJ-JV)ZXRDD 
@ JB5!E1 M50.^3377]HE:?C*%*-)2&3"EM+#T!8[I^< 
@;?/Y319G_BC?=A=S2X$\*F=O2J Q,4\X9B,.^'1ZF$X 
@0IZ8B$&F*P[)C=@];#$'\XBJ-PP$E=V7WV]/\0T/FXD 
@,'51P4M[W[<*]AM%>#8CCHV=N3U5=Z$@8AKBO]3OFO$ 
@%). <PC2A:% 1V(.?%EWW1K,7P:/1._P D'8.EL%X-@ 
@+'>^//J.[6[9BS4)&[=/0A83Q>\@/H)- \\S;M!"'"< 
@CK"&4_$N%-[8P0DDJ.DD\"GD(WIEP-8TV1 J+WVEUAL 
@_F%DJ\O,7_-A*=715.WA04IHW"KK!JY(S6Q_W"9C<60 
@[XBEY8^W+8:&ZEGA@9\&TVZI(O=5IXI'-7_G",K8O9X 
@#5[:A\8<;M.C/N"@DB83;?[<='?"@<D=!O7SQ[8A_$P 
@(L$!MY9A$2P;0^N.IS3IV);=HOBFO=X6_Y<OP6D]@ T 
@"ATID1.ELU;/]O GBU=5]><]_;=H[=:Y<Y8XJF'<CR@ 
@B3MPRF#II51:?] ^IOMR N&=?"LE25]42O6(UO]E^XT 
@Q (EK" ZZ6G9@&&^#;=:F)7/DKX?['8#A!I"13U@*/P 
@2A>F6P=*7/$ )]/@04VQ18XZ6MW2Z,1_7-)%4HHH5<D 
@L3T!3@&E+AR_KJ8+M[DM][AS$AX^#>GT[V'PZA/B1WT 
@(>SS@L[5#X!]FG#O,PDNC:BQ_8=JUG9X)<B'E=NBCE8 
@#R%^$NV&CKC-NA<E51.P1!>_LZ,N4LVW3GS3KQ^;&J0 
@@'_%#>85/HKEEYX\#!3P0>9?+7WZIF&21U:^:$SE%^, 
@HZ1S4GH*G3W]YUZ&C?HZ0UY?P6^2@,[0-F\NZ9;YUF8 
@ZP?T.?R-:]1L!VM4M?CS\]J6UR.CC9SR9+W"%GA";58 
@70IL %J>7%*=@&-D#5S_O1$*=CI,VE0'LZ\Z69K)=RT 
@<'SN7_!0:/:2?0,)^:.<RT:OU1MOLS49W8>%F\J^?_$ 
@I A-QR$AC%==OSL][UU5IDJ!5Z1E5>M\4RQW" D1 ,8 
@'-/7"IP(/=SR1L).(TI(:6CK@=1;3#VVD+=_GUTIU%( 
@MV@^91N(O\<0;L[H?8<D-:48'PX3GQ3+[N810SK\HY$ 
@4I(3(_<3J/HWA:K'B**<F%<D\[X(0U59$"RCR6C<(*H 
@Y@..V;]P9S^0:GY<$3Q'$9R62K4%],''I.;-="_P)J0 
@^*I5Q"?O$$48*8K)D3Q($77-\E*=L\1KL3V,6#/G:F  
@EJK+W#FXVL;V@;NU4=3!A/VO[Z/%<1R(6EBOH6>8-WP 
@V;Q6TI4QJJHT4LM:U'^R'\93BBL J&35J"4/7ED<=1T 
@M:=3-8BY-(WW2VH]H^2-*;4(>Q_O;BPL3>3#V0WI@:X 
@N@"B/AB[H4-K##F0WRC,!,R:L('!$':#>,7+5?47,LL 
@?9+[>+,R\Y>W835<=B+K6 ?$M@C8\"GF9F^Q269O+/4 
@T"#73P[;^<^9R6ZCJ+XD(C$:. K1*1=GF,L&KR25XW, 
@4>VX/:05*47('+NRWJ6IQ4*&U"J+C2O_LC?#!,%3GE4 
@]O%-':%#>/_&T+7/+>>%88 WFXR*NZ:JNZL?T%)@M)L 
@#"K%HS4\<'H>>)5FV]MHW=X^26M?^31_>BN+W[/>1_8 
@M0(J*>D5&B>X+769</<@!"MB64%CI BI6-MWPT^HSZL 
@DGUTIO^I4^@=SLH*6$"YZ_JB-<)LAW42AS^C3X,"&H8 
@II\$,8+C[-/%T.P^"$NZX3("._*KKCG5N!,@D>=^]]\ 
@/G&9=&*^['9.6Z":*Z-GX\D82@"PSM[$#M.3D<ALF^  
@KQZVL4]JX9UPI**]%$)Z2$_M_RH^M3#]+0]YIS4.2AP 
@@%#P!\IZVOS[JYEMRQUT$6S9RX6_U[,P8BC_9'ZQ4(X 
@= M,F" C?=:KR"@"H\!$'AV4@,4=^"Q9P_:XH-.33#T 
@J0P\ITI8'C!B7DSFT-IR. ]N$4[NY(6@88!\P0$B.C0 
@<51W!\E&B%?7=RO@2=<1)Z#XP?Z+\_[1 ^7(AAEM +P 
@/^SO?$ZN-ET\'-7PT'$RX+?X(4SXM+UK2)_ D9PL+\4 
@1F MYR6-"W)SQ5UG^'?+ 7G2&B#HKV/\V9CHI=5;"+8 
@ 0GZLN !,^8-U&3N9? :*@J)6,5 B  R_/Z2@R>/4&< 
@.''O$R$^:-L&7-PC%?YJK>4+ <;2%!B"1N3)63M9@\D 
@)X=3\.,499A5FF(Z'WY9C(U-^OA&65QQ9,,1 9J^IJL 
@Q=;"HC['GX!W7$2TWNUC8-=Q*[-PRCY$^$8CEXK*)Q8 
@LHL7TGUQ4'SJ$9^/XF(A 4#3+ZTLM?ST81U+;0NDSA, 
@S)Q#U2VGM16BL,<EUAB_\]_A RP-</_+[?PHH7@O.]$ 
@X9596F[X@+W.UF+$CP[,7P_2LZ6.]DM:$E"C(@,/O$$ 
@_O:M%=H^*#_L1_]7 S : M9'9=Q5'@Q1;)8= $0SPYX 
@:O.@(RAT;Y>G=&!!J0-U$(HT;'KX7*2: T7B(92O,.D 
@,M]!N+9&SK<<;P>!;=K6WJ#J/)).ZWY.[9H7)2QI@S8 
@SI?J7\1^B3O:$V0&^DM!-WQD*:FI(6]8C)85U@^7U3P 
@07WE,N#PH1,"\BQ.^]*;ZN,]HB>R6@VH'5(5$H_BD+H 
@8 S>O5\5UY7H!RTK0E,DV<7/#=A;%AI-(M.ZQ$M_9W< 
@;N)&Y]T2SH2N1WH\0])*B/V>*=$W;&U>_4+8"K%M@*( 
@Q7#U G4D1GS0MZ'9Z%%R7DS(B+4 !I%@8/,LX9W/E+\ 
@D'M-R[GQ2\['>3T<=,1O1;;$C='.Q46$CQA9ZH'W6[8 
@ZL%FEFRXM[9/[%_1>9!</IOAOV*'J>K7!*"PIN-DCKX 
@;8>30[._WAJ BD,3['_8DTE)W&+/O@'P$EIOQ?OQ9\0 
@U)\F6UOI!\BV-5/#BR>HO[2<3:"$_2.- [AHWH)DQ*8 
@G$1*LL6#.!MEBXI2"#-)%&CA]'EKMKC2L,*?@]+VEYL 
@D\UV)\^.[F4/1O*Z79::K1CO=F5K\ _Y'6] UD2;NT, 
@DO\)0<((E\^DF"=27/1YHD0EK(#?(K15>:,<9+&3#F4 
@["L2T?2T4ZFA_'[WSR3<$-!I:/VW[TJ0IP%?#C&MPA\ 
@+L-N@LE;KYMSP%_40*).4MO%GS>=O"<Q/:@KY\OK[_$ 
@[*:6Z O)RQ+9DE,_VW<T=9(4]U35D%O! ;GLR@^LFQ@ 
@%KO[>R(3DS7$+,(+)R*V$K+:;HZSF=QF_!])_U0-:1D 
@&YK-*;G#J\>$AIQX5OE:1-]U/6"FRAS)QRB[_81-IP4 
@2;8L>>WK.B,CO<NW,F;$F79"G-#;>4A1IMELTVH70<P 
@PSL45\Y@H!O[%+CC,#>Z165NQ&S!&%'2YO7EDE!!&;L 
@..XJ=16S#Y 0I;SP '(;ECY],VS60.(AX%MV+:#8(0( 
@#\?^_>D1R>0P0SJC0V&!R7L?7LH\HP]RW&@$BH]W?-  
@!='"7GSR=?V.Y-V2(H+9"M-/ GX5NX[A4#;HIL,47[( 
@U+F;02TCBIDLQI)[SU*+X9 3^%Z1C2&%8"<$XZZC8UP 
@HR X1#S=L4>\[E'[I("G\ *'^P9Y5SMWV8]&CLLU=6T 
@=+M4:\3 $<-TO*I1@$DQ)'O8;;$SAW>S>WBGD=Z46U8 
@H7K(Q4M#&S*SPF?92**T%)-S(!)8D>>S%8=FY/F\NTL 
@"3P3#+B/8I/047W\[Q6 6GDS*SD1.1[N6R6@=K!$ :, 
@^3]%U;:[EV_ 7C[Y<<#%&?>-/5V&/4;)9!]B]<XLC4L 
@*(:I*BRQ=F^1ZEUEI2/*7RD*!^0.DHW%4A*]==M3%40 
@C*=S6L\?KN<NIIUD,HS7I&B.\S_+D"0O@L=/=\993?, 
@@/BBFI+P+JZGQ%IBV5/^,L#@/F=TLLW_HN>L"/,7SD, 
@K!-939]FZH?Z)A492AI*\?76K<BCHRQT.B]YP-[K[UD 
@I.%Q8[N[]H]"G67OW;=?>1QR&F:ZH.;#RSLG^>MP1NP 
@.6&?H\"[?VO/-$60\SG5\P,R&9&1&;&@LC=\-NT73>H 
@^@#T%F2L&'372ROWVT_B+[Z#@:6EZCZYAR+@-LH1Y>T 
@^_+RP L1.6SHW^1AV=$/WUMY^$M?:\M9SJH2'K(N;^$ 
@".%H*4Z^;5B_C"J,/FM=*F]95O%E$+6JW7J([]#C>QP 
@<L]6WZO/2IKA_J('"S@F;6#G3HWP!52X?TUZ<VN(P/< 
@B0?+QT6!UWS?WZ]!NW$];RO^^, 1#045?^&NE-:_31D 
@(3,J*S?!1JI37+\UA9;+P<)7PLD,C(IWF&0M''A59 $ 
@\%/LG7:*+BS>"5LIT'#Q^T3%S/UJ4MF>,83 (T:F/V@ 
@"_<<2G8EWUHUY[]/1D&^YXD>T" @('YB6#3;Y%= 9[< 
@-Y(.327:O;$/HAH8<F?ZTFC:_<>"'@5@,)F+DGPS)TD 
@33G8T%\4.ATJ9E0=VZP?88B75 M7N<9@#.:=("&W\<8 
@)GK1A[D%W\QM_5/6/KWKML_TGM9 \M)]"U'**/>"Z'@ 
@<!/%ET_*LN.G_WQOO?]X E$ [NNO[<V"A@,)^B+SV]T 
@E!ZS]8/QH_&[C-?.]UD0ST6=< ?K+U4]^OA5[H_CPQX 
@:+@A";>T^BR$9G09IH$P2QQBYJS-W>Q@@ [B2;0Q!R@ 
@5/?$78\2,OG&ZB\AB89LW+!1>R#TW_+$)UDU=JXFC[8 
@%\G9_1-[.XD8-G6TX;/C7.-G,8E2L-BL'>EX"QJKED0 
@P&%+.'9)!MIPUU<<L@_&PP&[]*8,F$CJQIX7,A$!;!P 
@RW5C,FQ:P?S1+B\X\,<?$,&#UN"1TH0(ZUD!U.63V1\ 
@A$UHD34(@]KQ\?9A*1P'*VY^*O,[L]-C?1JGRF8[_<D 
@C).I[3/F6_\@(.4O3DSL7D[L)3$;([0C!VXQ-SRG:H, 
@Y4%"99KV-\N4W6^AJJ\^60B.UH"B '6[=9Z+-LX';@T 
@Z.\MJMA'%[$@@>;%/OW%53 5N:Q;*U(FF/+[VX5L$<< 
@=C/^];@5(UVQEZ8*(>V9W%7)+BG:7<L2[3J[VP@T#O< 
@GJ8/WRM6'TF-<)L.[II,0$*Z)JS]46URSXM3A[LSU < 
@-X VI'@S&&%#Z8IPSF>+5#B$GA.#Z$;UJ'7_;*!=J1H 
@4/<[$BQ.B %O0$>&H43XAMO^2T,^RP"C. Z6/8%NLD4 
@@=7(1U3Y\?6MXH!3G4XHL;M[8>6/ZK5]FNQ7UE"DK(0 
@[;JDTI])42?UD6Q;?V? T$\S_ONA7,IWZM?<+ZL^CJ8 
@*#V?X(*IM<M H;\S,V,9[FU)@F8C&J$'NYQPSYJ+_H\ 
@=,2#JN=BKND&5U Y^L@FU?AT7FG%*-4N'9?<VJ544$\ 
@Y.^VLY-[K18$>2U(6T_9>M),U2W6VB=+N,*+6R#4'L4 
@@&XH@OT4;1>T_U%H.<Z1Q39PID64^]:E?$VX@OH1.OT 
@]BC6=[D>4Q;.A\_\[&<(D" K^K:9&9H>DB@K^;7(VQH 
@1E6X7?ZK</(;I4+_U4L)DS3$DSH5;2#FHZO6KP5VQNH 
@!TN7*)#Q%;@2VNVS"&RT@?W2.M2"1*+'4X;VU1GQ2-0 
@G2O/8_;7;_98>/*=U\LL<=)8#8T#H(6@GOA[!GB+T 4 
@O3 >]X$1'I844^UK-+8EK9>,LM8#PZ%A9G@BA]<X?C4 
@I +M31DT"#&&+?>W-PV:MYJTU:)H'FF'QA6MPRIYKH@ 
@=/0PARE6P),\]DM?3S[(M#KJ_%Y$I&D#(N!2Q+PH@/  
@4;QBEVSS:@<GG[F)7]$8_[^2ZS !\/W EWWK#Y/!K'< 
@1WZTEL>0A;!"=E@-]CC.*$_]E!P,]=O4C3D,W;EIVKL 
@J-E<P:_$,7WV R(9[%!'\PFBBZ6AD$$L*@]+]I45<I$ 
@#=J/7:'P-6; *"$Z%RB94Z-^1"#E+SN63#8QX9#8$D8 
@@^/0-BR]"L#$%GLW+#/8LJ6?:ME4$<O8<$CN'7=,<-8 
@T:6O7VQ(Q!F5P6JD0TW7)T,GB,"D(A2C:5MU!>?$X"  
@17JC'></=PUSZJ;W+JL#C":<DN#MX'"W#Y+DAN+R"7( 
@.Q-@%\O)%@H8->][<LMN1@%>1=N3F:ZO.2Y)*K<:7FX 
@%LS^DU+5^"M1>:)Q^Q@[Q"KI5?TNK&^AU-+*$$EA"-@ 
@$U1)+X?:=UGE0B=I9NR"V;K4LY10C:3FQ?5X.Z,0K0X 
@:\!:G"*3C51*S'PAP?5M;!X!VK7&208<I8]1D9?I<N( 
@2<#8/AJ(#Y0\"?,XU>?LP'H1SLG!8 4S$H&*SL]V.X, 
@\ UTLG4CEHNL%MHHO$^:(W!Y&JX/[C8CZ:I<]'7)B<L 
@J _#(7F(-FI%R.NIJQKUR3Z]4;3Z=&S](O=!^\Z!=[H 
@A- L?;@71I^#S<&+SQ:TT4R> !(XQ>LN\JL+C=)$F\4 
@&ITQ4U4Y/18:?'()SX\^-JJ3N2=8KH5[?C"YPX,&)XP 
@;,>[]O:?(>CG51DZE0IGH'@ !&;AO%-JF;R_3=R*]I8 
@IW9>0!//$MXRD3&VHCMS"X*> ^U0N"V?&%NQ8<3\:?< 
@@'D8+P/=&,#?CXFC4CC,>OA[>_C$_U\$UDYQ3$XP\=, 
@9=YQJTL%0ON/G-[Y+5HJ523U;&)RX^@$*O!\]%&D*3< 
@;[U!@+]$PE02(8S&VB22@5&87ZV5Z9!RIUL3.W\6;8, 
@]R0N+^>,NM=@U]KR3NI'UKP_'X0#T/R<K6"QY!G].@4 
@A"]DLM\'7"G?$.Z#,(S\:MJD#P6+ RM#N=_'TV]EAH4 
@P4Q\''WK1F8.7<7_GTC4;_?E8TP>1\)3A;X<GV4M<<< 
@&%YE5 W+W27Q%7":DPIP;XK(N->MDUP147=UF/';P8P 
@];@?$(?5++?\?]>_BNJI,_#T!^'2!UR%EO"ZI_[SX\D 
@>!LDD:L"H52PF<H,U#\.*.<G+]S("0W'C5;P\O/#S1D 
@ "ORCJL:4R<189IZU+T*SY3-\^DA5C6Z644ZB-HL'!P 
@XG)26RA]>V"K8MY?MI!=[( 9(OT< _4;]T17ERZ^@ T 
@G?6NV2M,.3@*_[B:1C!0R.!Q'WTV%&YP1[ARY?:STIH 
@8X5:&;A[0Z?)\?=4-((SY*\;-)6[RH#WOW$NB/BRL_$ 
@0+^#B\E\DX]R4G7JN+#(&H83\1YC ?@,07:W9QYAY_X 
@/?NJ7L'KW=]8/K2H]RSG*-1VBK,BW7S [$OK^;NJ* ( 
@S^-,P)Q.C]>14PXN15@^;GSF+IG0P,5.NEWN'A&?B*  
@ [UP7\*+K8J1T3Z.T.S?JRRYX!FOIF=U1O6>ASSQ^DD 
@[) 1T,OZ>M?M5&U W*%_LU98HY3AJ6%/X-<\C\))4*L 
@Z\H8WO<[0'3@]"]CB8S\6#)!"D#_CYOL@NO"+B(Q;], 
@R/<+I-2Y30H'X.^:Q>-@1<[O*,<78B/5 J7_8[ZJJAP 
@)%+QCW&[9!Y($16%89-Y_ _A9S/ T;QGTJ%!YJ,L<_( 
@#A'Z^G]B>IJB;#R\8AN6/<<OZ(O_ZL9'1-\EGFFYEE, 
@YDU92Q 1=WQ64QZ5CHGU>3W.R[@GE@A:=LBSW5VT^:< 
@15E)ZNB=&1F/JQXUYA"\)0?KNZ4R<-I.:F34TXC:MBX 
@JUK\S&@_4[H%+[KM,KJ\Y]0OXO"#Z5VY@6A\$E@T\$  
@ W[#E/W?YXBD^Q?ED,'K(.VG-:G*#OOAG>59U@\P>=8 
@30$+(%CG '59;6WH<V[**"*))+7HP4,5T]V@GHI*<#@ 
@WK0PN4;1&H?='>_-TL_!.Q?R&K.7G061K]>UMO,(E^$ 
@ML*5GZCH&#[0<FMG,E=.V2#"4YW#4DI/</_]F64_\^L 
@L'J";]"NA_VSE1G;7F7#H!8R"UE]]LT6/K15<0>I^>0 
@4%\SR!GRUZWZ1 0]5/M6GA0(Z7]R'7OBLH3C4^^QQ,P 
@-M<Z*,\I#H2 %RJ$=4U5GO4J?#I@=8OJ1NOG:^\MA0L 
@V65ZE\2B.?]9+&]06)D#"4#$$!7$X.+;<UE'6CQZO(H 
@:M'L(O#/W2978C F*E^K_^32US?#UT]4A]:'3LVY=%X 
@L!;^:4YVD[-OYJ(H&]?2ILF4Q'Z\&L7?-D8?##5LL7, 
@/5F : *B)C_'6F[IM,.O2Z2[ ARXH,+V\(Y].S]/",4 
@7XVFR/W?();PU^N#>PK%<^P,@:X*S-['3M[>.#W5:;0 
@61TUT]QV\Z%/GV'M=^_EZ:$&*%BED:%; E^58Q-AG=X 
@0OA&6QQ#$Y9 JMU"3<4//D3"E3#)Y<;[L8CD1MK<(YT 
@7IZL98[W0S0YR7?:W-V+8H*C&7H>OG)PBFRZ'MKTUPT 
@#8]./GY)*0=R=X0.@ZY,#>!;8&AG;-T:GLO,'=NLRE8 
@%12,/-M3O S+1V8^U$XO]]^P$9AXH[MQB?OIJ/]6<=< 
@$=#*<9$)2KA-.5NK=A;/&5)<(F_A=NE-8]?@UK^(-S$ 
@A<:]N=0(W7!SB#6C,)AL/?!I:^LA*MB B>+S^D#$S&P 
@JEH[ETF#>]TTN6K7DEJ@;0ALYE@,>6%439<B1M,4NVP 
@YTSWX;BG+C/6JTI*>:(4BV2QG4SF&SHJ]L-?+I*4V^0 
@FO=,S2#]:6F\+E'QLDEI543-TLO"A**^N\\4@\!IEBL 
@LQ!)[$DW&]+DN-C1;QZD%=0=-W8M:*N0Y$,]@Y/UTHD 
@+]/QU9 %A*^*<Y9Z381LPPLMHC<Y)>HL#_MW?&5&'=  
@N,X@D\>=A#-16/#2T4U=;BM C(2 \>R$5%YQ\'90[!D 
@B<OHG"3U!&WOBP+9-VP?N!T59*%RXG6@U&_.AL.3A3, 
@MSD@EY7G_:#A(N!YOURT;=+ND7+6U>(DY0[&+I)UZ#$ 
@2=EBX#&\<: D7H/0#1&E/OHOGP10%9Y.\7#MW.]J,&@ 
@TVFEKIZQ@!0]=,B>*\'69-A%](+%+]#4@Y2 4RK""@L 
@>;2Q/H7BC"_W ZZ\Y )E;QJ%-)RN]R!4 E[YPG!:\)< 
@PDW5R+MK8[=%0AS!XM.X;.:I(IG<2 ,Z%/0%6=LY]I4 
@* "D5A&UAX@.@XD(OHD?M)Z TQ>;]NKO'[9MRL*N8*0 
@U5TP].BIGVQ#Q,KN^>8L1M?4X5H\STB^RLL\AQA5QS  
@<4*& + J4)_9"[\2U[S3B?7*QY](;D)D<^ZH!!*'N@T 
@4@9\.F47Z]7;6T@[1HZ[NY48@U=G9KY9![!2^3NU:>P 
@^O+0KCN']P[.W<SWP=YQDUT83LO+E2@.P1)@]3_/.;\ 
@J>22:@72=_^#KLA_=>%8V)OJ]>(S5BYX@#Z-*8);7$@ 
@@J)Q M,.-/GWRN??9W/_(YB.Z&57RX(ZPNL]#!W$9"0 
@62,1UZ%R*W%6M>CDGVEGNIRPC"2E[.!0S89)6NLY>UP 
@^K=1*/$D]JOM$CXBA(%[$5OMJ)=W2J3N#?1JPK>O%\, 
@V9G&I[X0G4. P>9COM"E&TJX>+%[U%.\"\]BT3?!R@H 
@_.@Y= XJL3'!%7I62#3K,*^&^B<V\O#9^K+"'VJ\G=D 
@849W3BB2EC=N?L^!5NW;Z3"4:]@-*>L&^E<P+=\!W10 
@11_[3ZAJI0>R(M40E:O0%E'. R=.BYH/N>Q)"V(^9AX 
@7=@XC5>)L>6[G?,Z_BV#U]K-: O$8@C9DN@L&"#/,44 
@P\PWX@B;&'7DU[@J XB@/X%_Y@#I'/25R6B+<!5OJ[X 
@PDSC 1\EQ6="K)"_V-3P><2T(-0 )9]&&V^X\NG>"4@ 
@,C9&CORD:"M3H_16*O50A;&0P(7N99RMF95?AX #+?$ 
@'PJ)ZX$=?\8;&.V9G)(6=H($#2;1VG@'2<-R;S8Y(/$ 
@G[M+TJXNH#Q)>B>P=LOF4J7V9W%*NLU_ _\O#%%?6L0 
@C-SG"DA6B1E*L^9)TN$!Z!X\*)AY.X[!"E.W14;-13  
@//4(RM6#OB%C/"M'7-$#V<41!=!?W@V^T04RF7K+AJ\ 
@']9SZ9\AP$NAS(";WA T<FXT];]'R#M%;+J50HQ"RX4 
@.C1UHCBJX70S.;@(_+0TD.N[/QWB(T6/'K<UEBY4<H, 
@_X\JZXIHF B$<D:'DQ&^Q@L(^1M%\W1_HY00-W3 /M@ 
@%&M3((?*;>3JY&@^7*FX[=-V0S(<TK@6O?MB9&S,N>L 
@#%=?%*E,*Y7;X8(=*8.Z#+;D-6#SH("UN)V&(^ML<E8 
@S*.$M]3'\**9/V<KAU]YLBU/V @MM5O"OJE=(1 0W,H 
@MD:+0A@LJCO*($$_JD*X6L=057@Q)740,M EKD8PI94 
@SZTMM!R)N-[6$U9L TO:RS*Y7QJ9Y'37X<E!#NK$!5D 
@AKE+3%A,GV1I/W\H*/;?MB[YL)37FB: J7;%*I#NN,, 
@+N>#@8*_]Y^9!5%J#/\?5&O@P%H+Z*UC452Q!\#[R)0 
@SI'V==9W2_(2K&K;W Q5]8?GZ7%\5]Q]R5)&ZC0N@YD 
@*.5'UDE1O,U?<\_B1+K:;_R^M=QKO[G0<?*'BGE=;@T 
@JXVS.[*O0=/>C$S&G[)RL",G$ED]="L(IA2WG?FN.^0 
@U%*("\Q%F;<B<Y%A_%05UBO$-&Y:A:U5&9A693/@G3( 
@'+\QH,<X-$$$)]/Q/>+:3Q^2\2>%B]W[E1TX&(CD@64 
@N_Q$ENCQJ$G/(NTS*$.0[4HE7KBKHB?\9I[UA):(#1T 
@C^]MH>1<GH"M(#;FM]\KZA;CNY*<?&-\AS3W?&UO>L, 
@YP.V+F*^)N_CYM/E%?#S2&L]IO"@\+1;='L/>"=GHS( 
@]CR )E@RK 4=\NB.K77R\BJ=];Y+)E07B\/\-:2%YD@ 
@ET" :%\R\?EI=LESF<.KXN2MH1%]'OWK& 4V2N;&? P 
@9_S?J?>:NCKU+&WGMOG)#P$[D0R(EC(-S:\2!C O:7@ 
@/#HSG[U&,'4IS(E4)R;-?HX(H3[(M44FK>;IMC$S6AX 
@[Z1BVZ*" ,A:2[XY3Y>7(G49D8[,$8IK,^+TO'<UU @ 
@ML^+S4S#+!!C+>_!)3RCXCBDWRT,G=P<O[E?Z"/K9R( 
@3\Y*$#+$G+9&VD6,0X+>3#,=D]DDYZ&-6K4Z!C9K\HH 
@AZ2@2GM7^?'B7PF^5"]2+TQ9!)OH_784^'R:]=X]DJP 
@_"+;SCC[#:L3/>-Q-H[OXB:#=]L$L-GX3(E"P!E (%0 
@E#C#7]/_<$W=W&RW, @B&B#=PU$N?#FT>AM&]3F([4( 
@+ ]:[:)VVY\33B@7F0Z8,I%Y5M %T+Q+Z^>_%6/<W04 
@DIVTG9P9+PFG&5_K\3]5!!O^7)@5S)*#UB2(N['?OR8 
@JTO@@8HB.V*J_\:S/_P60ON(A\YNSY'X,W#YD1E9<[D 
@9C]427S04G%(9*^]=]6U%YR6-5ARD(@$HURTM?KX,=H 
@U* +\(?<6%T%@JKU/2F5]]Q ,4=^Q_#R3I1K]_S&<S0 
@!$W<J)@M&&MP<3@S_%S"[HMWO2)7M646=%FJJYY"Q $ 
@0T-;KQQY-B@D0O2-!CT.$EVK+$#WBKS8K'">HRV3' P 
@?0"8/A*35=3(XS+3ZR.@)ZU7NB&UQ'@=64S2M$.T<8H 
@CSO6(?BU5%N&OGK(4C^&0<)L&PQ^$7RVTR07'>0C4<H 
@2K<X\JIT&@.\D,HC4W\ M;?>M6[V]CCT;K1 X:&F:<< 
@"V=!GUR(!^./VZ55UC#OEH2LIM!P=,,_O".2/^^O>6$ 
@*66?(809BA\AQK$FD>!4@&9O#9#L7+\G_-X2@KJ2D7  
@&=R9M/Y#(1S\X]#U(QD4[^$*T+7@7X+>O-53<2#@\TH 
@57VA>8DG&*FC98K=3]=@-WP"]2*[]CNN 6 / 3G8L6X 
@/(! ]==U![HEBFNA)KT'A7(1Z(+1652U_T9B3NQ#*E4 
@R'0M]4F')L*[_%R*T>[;]/%40"0PFF1[FXDC'CS;2S@ 
@(3^UPR58*_MZ5;UTCLULK$=?//^I_\SEI/HA-R5:R"$ 
@IXMVH8I5$44@ UDQSTK;!\9M3G:PR!F4D\OQ,HBZ&30 
@\6E1@Q;D8RG-NF#_NM1<2$A'7L0^1<2C1[:V'6)Z$+< 
@DP1HS4D*G>P/WP5OP8F:=0_Z8FEOJJL!P!??298MD5T 
@E7$;E6(6RR3KDHJFN5;?:\&T[\MNF%/TST]8U':8'C$ 
@F>)V7WD'V,[W@#L*?^.7R^1K7+M=F (WY39FY^(?OF8 
@)+7RC=!U&9%!RY]QF:=6^KV_DN,P6_8[F-WN.^^F]F< 
@HN&J=R]<;@%0!+)O0%,O%[WM2^$KH[^8W+7YX>SM<KD 
@B Q/C&>O=QHO>[&(&9P' _"I,7]5XXP:#:WC$2.?9^< 
@[\,-"MM_:%H(-Z<RBEL/=@8]DM/\&G95 >:FH2XE],$ 
@2RB4G .?FWD2WJTC&&MD@7CX?'08DQ;4X_FQ+0?CZL$ 
@<C=K4JL2"9W9VM_P*^6!:=S-JFJ18IT&)18*QML5AK, 
@Z9N3OXI1 I"A0_F;;F8.<$T@K <MB4L9$$-K44\;/'0 
@ 1D8IJ2T7R"S[?]5':PW3Z+I^$I/M?2@K@ICS+X;DP8 
@!.B0 H5B&:!8CP.)B?_N2=;S1X7XD59'BQMXBC#I:C\ 
@U*,Z(_!58MMHV_5:(F5:%IG,>O_L60Q61<Q;H[[G2O8 
@7YD* %E0JLG-P;E*& 4_9<:RU9::/+F>B,Q*BQPF7"\ 
@9J$R^S*3A;!%5U,MKJ9:5[L)+FX+]&IHY:9>>[W$IH  
@I#68=V9GB9/CD#$6_YP&%^]]?F$Q_6M]W$#RM /X+@  
@(_^:9%^MRFXU)$TYM@,V4+H&Q=MN1CC=1YK;HKM4\F  
@TI=H! OQK@E#/;'CDLK#8OP@RS&G]L"W!:.$YX5'X(D 
@5#Y> IA-#E=)]M#DA:1@DA>T_VG)U;##^'/,A4:_V9( 
@XE21(1-D))[>O5P:9"3WMYQMF>3IS' A_OD8!%<NY0$ 
@OV"N@.MO1I.OC?NY*SNS";Z#<)01J(K;\SS2GBQ'K28 
@R::0584*U!"MYZ"GK>NE"1I1CGI6YD.R[Q&*8>&.VL  
@D",[]A'/:7&+ R<FA<N]P2<"".S*5+_I@6+LIBR,@7D 
@PX(UL0A#.>)W0U>0*/QJ/0/$(0U%$;A0"_'55-YFC!X 
@.;@6Q=ZE3-_]]F2DTD$3CNKB'4[E50)^H;9)#4@<T-  
@-8V-LECFG0]YZ[E<6*B5JA)#078=%^$*O!MKOQILLS< 
@AO]H3-<IR>32[1!DQ;0[GSN@,''8 T"5]V3ORM8C@ZD 
@_Q6GT^?E884+E_//*B 9VUZ!P!9>YG4LM4N-H GY#VX 
@CT$L2+9_1Y:8Y*[1#,M$V3.Y@QPWX'BM9K<]?E\N+CL 
@SIY\@CZFX_#W3I!=GH&E(YZ1(-GUGV"%OSXDDI'#F(4 
@"3&^7GFABQ[X 5J^^SA@\A&U4PP2W<5RX"ZHC#>(:Z  
@]]!,EL&?]/*":8PF99(=Z YIA0A3O1T*X3["8"_SPSL 
@<#R9W$_V.F,O 8IX_+@+#(__]#_+!$A3FO_RA;0OO@T 
@>9MYVEB/)!8S*Z-W#6;BEF'-ZPUB#W,BRQHR?S)3&U8 
@+0ER52T%[2.[LQH6GY3_&G=_*>6!?M@^6L%Q"%W*_Y< 
@=-CR@QT!),OT,G-N;+BA6W3J<>3$1N  6%I127P$OF$ 
@ZJ1^R=04?BQ4B1R40^D^7#J&6T+[*BTBKPCU6L1GYR( 
@";V9/.C!C>WDPT'_JCEX@1:((C"1&38KS=A[JN.2\:@ 
@ "8%ZZJW2?FP7B0PP#J%9005[(VJG%'2SX@2+N)DQ)\ 
@,E4#5"-  *]<0E$D&.,/$])TXM^=W>701-<*6<H53PL 
@/X:F4"18[KH%&ZB:\QS0&B_E'=2+J7KOC+?%W58C;*@ 
@QSCZ<VTL=A.G6T@.>XE6@B@<HE%_>%W_*Z;=Q0GSVY< 
@[9B:/UGA.XSA]=MOK'S\SDDE7C@H;];][2WNX1P%;7\ 
@359JG_&';MZ8#P+@@6,GFA>!IK'KW\#%C0OE2,;^W!( 
@;78%I(HME32Q.0_V-,5G+2Q;8\60ST)A>%;00FU7Y2$ 
@8VF[Z4F5K6,$J$9B+JQ6CU:E]PU?JENI-^W\3^T*UBL 
@VT,%\^=G-*WU@<7K40;I3^(5&T703&:[?188*%*@R?H 
@BD4AC7*M+1A/ZHC_F$X7Y&NSL077!D596*'<<^,<2$@ 
@EZ[$9$38L4_)VBJUZ;9Z0;XZ%'/)S \'*/I:MW;]GLX 
@92DZJH/V -DK4XN,F([KF3IZXLP3D.*Y ^%X>_L;^?$ 
@X>:<.S3\\MK\'&!H%43&D6<FR^R()"\@Y:M/OH)T?80 
@ :&'77^6%^4*47G]%V/3T_;DZ<&-"X?#3024$B'?N_  
@\X/TOX%=-'-Y]"PZ?IF2A(@VV6LC:_;SL@^*277C?2L 
@?QZ4OZXQ'3W8]] FI%LAH9CE+#XNX@-F.M:"B$;033  
@ +6[8X=Q[P] /J1P?ZFD(C/8TV5(M,V$94=5RPTRR#0 
@@F*7<3507'=G4J==305H#J03W*+&R&W@ZS4@SRJ^?/4 
@WOR<(V^(V; O1[O[_V[(3-;@0;&LI \9L_T7(?OVB$\ 
@GE)@V=75F+>MT/@XU_(.;6IG@*NB<YE#E!0(YO!,F>P 
@JK9.]<ZQ^*@0&:0?UAHPF-EMU&Z7[?D%W3SVB'L/+DL 
@3.9J8ZEOKP%2Q%OFE%8@8O3OZ/>$]B4$KB.2<\ M_/, 
@T5"K2+K\?+FJ)SQ[;I+V5*N9%*XI3?**T $+;S;'<!0 
@=J\,USW 5(4P)'] -SQ SS(D:<?\^H/@_>=S=N:9#1\ 
@@N"@*:"=)MWDONT BK='*%_\YS]=5504*3 0&<FM<!\ 
@%A,[VB&$&\2P7#F_UP<0SZ-_R(B'+R"DW1$%#J/*U(\ 
@CR656I4,WAKW?#/ P/Q$;#<_<HI! 5 AT]J XPA$/B  
@XR7UB702F+BKGZ5PH[OY909@'MSW<(L..(@NLG<>M^$ 
@J$7 X%M 2M0A= )FB;XW<.,NRC("7H]P?O8K">PY+S( 
@$&5&CUGBJ!GBZJJ54TQVN%8^<MP]8<XP-@J5G1^TC%8 
@C^3SYZ Z^4\=*W?F#"68LOM2Q,M%5RF6:>"5FZ<074  
@\?$K&*2+/,H(^6KE9!==!:CJB9S!@T!PHLNHU)!K3EP 
@FK\'!]Q([5Z'" YZS-G?2A!7C-(\9')"3WT@.T3E1FT 
@E3[AOKXNP#YM2]_?<C&B0@S1I#7)X("ZLYYFJ +(1Z4 
@(S*H+IC'LK-CRM2X+RD0O@%/B,YR\VLA4JL.N<;5D10 
@_</S/B9E)D_RV.?:D:PO]N@Y$^O)@9233VAR5WC?^ @ 
@+IF.Z-&&P9(FS6XFC(B#Q<SR1(W[Q_Y@K+H@79P!=7H 
@QV.4$.B<=:[R7G?3!;L.0^)!M!!,>+!YS^4 E;T*$&H 
@%5BCS=7W 7?6:66HD H/9T!MH3G+ ,)8)L?H,;?/ 7@ 
@NQ_(7>'_\A@+8>IL@GSPN(/COA[TU@.1M-:?K(,8KCP 
@.++4MV&.B_9A!W$P>^: 6/L+2.%89,MV1-"2NLS_9HD 
@-HS%]G?#)5R+OT'\"#M].+L-..@,NIN1<,T[X;1L\P( 
@C0'(&ZC.Z^W>$<;WV/!5'.F=PPNL>Y.VS8U&#O/12 < 
@(@95XK!L3U;PGG0PB.SJM'-$%>\>"RZF4B]LIHA*.I( 
@?=\0(+@0C/!7.8R#+QI8,YE'/410:S7KJ0XR)%VP=LL 
@77AH.R(LC#1'Z7]VF];UK?;@=W<6W,FE5F9Z-JAB.LX 
@JQQI %\!XB%O0ZLMD-99W$EF"QE7$.+]FS\&LV16EOD 
@^ I]^D@S8K6MT2?1JG8S<%"IH_^L><W(.X/G" DSGR( 
@,B)EC%>"H>?,SU),ZT*?2RMY7EC$M8%P8J=1H020EK, 
@+C@.SB;O=@?0=_40+0HZ6'I^+!=7OFY3XQS_KM'^Z40 
@9+:1[>LG>AK(PR: 6=QX-@D:MR8?;-W<#;%5EZO6#$H 
@69Y/I6"YEW@='7UU-,X_/Y?\A&!,X)3&(%/T1)_?'B< 
@LX[RUC9X#CSR]A4S8-4\'[#=[=X=283)D<?JC(\7,HD 
@;A/V>?$86SD[I$0TZ-$IAVMK73M=$UBFT.NJG<F<8E0 
@[SM(:\K)^Q](!0-@7%N#7L]_MO!@-+=G*G--D:*N*#8 
@QCQ[9FXTCA08T"J1XA8L/B#F?P3VHT9"V8%TA(P6_.( 
@NWJ?67\IY+\03S.4<TM,3=R!NFMK".'8"W8D@Z?6=9, 
@BTU>3Q4#;MU4]I?5$7A/1K;,9^6ZZQ_BH@M'^/9^BR8 
@&@L?'-EF@1<@(:3.B\>-41IB6::K=&?JO(#7% (2U2X 
@7\IH<AFNY18T$EP>J"9WO+ $7QJ+.QWVO 6;Y@M&FB0 
@@1>0NR-KYL0S);GY.EZ(K(+.%YQHK'>[D;.ONTV!F?\ 
@A-\!J.WU2-N=<4A.QQC7#F- :@QEV>2<B@M>JBDCEM  
@OYJ3,DG?H15+?V:D;*ZU>*)L\?4M7)^>YZ7^DVH=XGH 
@4[FTN=;:G3P">[V9ZWF49Y<PF0B^<)TN%FQ3,;CQ%!0 
@E;*R>WK'66JI3^K *#9D)-"#L?=ONY"%-THM/P?OBG( 
@#\X3CE#',I[-"'W.!;28O>5NIDIHJA.5:%H-)=!+OYX 
@@*H+CQ1KBK7_.(WQQ1?_=B':_\><F7 1!.1]PZ\<%G8 
@>T[M>5SXE484=L BL>)PL.^X@ W9%_!AQ>;7A/&#PX< 
@+$2 4*9V,O!U"];T8I2*)A83\TK FYI&0ECW<K204EX 
@Z?"@<YQ*D3*DHFHD 8ZF/=I/EYHUTC_OAV& M:]VI@$ 
@4X8O!-5[;(T_13MLN$PN+$:NN^2$!</X/TS<94MU;LL 
@V1MVE?9@;[FR@\'S^]UK?/D]\KS4JFB0^.3$BP6C_EH 
@-R=B= G[@HCR<*5VE#C;OC6M\/M#.ZS< JACK:4/H8@ 
@#ZY(S EN6V@L6 ^GD(>]TSB9#@77<P./54$O [[B2N( 
@'$COI(+)K1D%#1KZR*;GNN@U+*VX*CN7^A]FV#.CH2  
@Q$#1/I_APJL;] #?\VA+M7U(]>',-B8TBSWC>N%A8N8 
@B+EU:FUP 85PU$-UL<*-LR@$#7?-B"JGG9HGAZ'=ONP 
@Y@?#5IV52@8MSD&"@2]L,7K/X%#SW'CG#V_T]63V/CL 
@:/]7)(%KA+Q/YA#/0V\7_XABQJ'<:I<6EO.-%6ZD@RP 
@IE@JD.,IB"H)F6]$C$7,+G'Q#[.)!]XZW>\&5OE2S!\ 
0%H&M78R3>FT]+;'H#<1I_P  
0>IB1C8;#=:U$U.D-G?FY%P  
`pragma protect end_protected
