-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
32xbcIk0+bL8J4EyDI9Ze9jV8EsZnoSSGjYciua4AQ7OsQhIkTEC0gi4iUnTc07l
I/g2rVr7Sbdv9GAEZbVEB0Kdewx77NB+mBSwrAxWX7GgVsbVM8SI6Q+rzZ9YeLX4
pQeoo8j4d3061dbWQDDh9ZL6R8zuYWdCZNk862LQd10=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5200)
`protect data_block
I56mrXXG8g09/EdlALYBBEdL4x62W7Ch5P5+LpfgcHB3JVQOIku3/8amiaJ3sICk
wOIHcQjO5HZWM/wkFKgUjn3/EcjwkjUTZKqVrZFGNwBY7/ZryjnzQso5/o3JWDs6
O2PtDYmvBGVjRJTjIXihc3cZSzGYtCtx+fRsUx0MdAIM9EauzgYthOYUbnL+pmac
knHFASscPCfxicwSKocN3Av9ahXquXKAyoN86pBywCGzKG2i6DIDVY1pyMX7ixuE
wLtKQjkG9N4CH6GU2FBrnaLbNtbzw24U4RJAzjobIA+px1MnHlMELtSsyqpqI5oB
amC/djac8hsMl/U4N+Q+d15wpIASfbOF6sSOClw8B9632MIk4NwjEZLS6MRhUaP+
ginwaC9MfMuSn7pU0VIVtc/UUSdQ5tjhCpaagTvSQ1q+tZuBXzqV4Tf4NgHXnRgZ
OoomwwWKYDf6icjoF5o/kGJtApp+E+L9ZScqSeSI2PXjCaADOVDkQ5gJobRwfyJD
PNknhPDSIyVn97kBI3ESOK/AeBAbb3m3aTwsrrZ29Jai3nQ0SDX1JXRhfzB20WMH
rZ2aFx6CwlxTmuiNudQOWHEhiSp8j8ziuZvOhVAEcbPVO/9ajopKnS9q0kBFYQlU
rGr81i/zir7P4oqiln6T9SLOuGVSWKAI3zlhqMVceMVW3f5aMLMFtvyJt4NPMKKl
fZydqAi4v84eR+A8xaK8vcaXBK/CIlHaai7XkLPig32ODHgKX3pHBTL899nfc33Y
i9a27JKowPofahMMfUM72XstfntCawyXtU7+4DvqievwN1DAYTOyjgiupx7t6TAI
z3+Pl8RzVBZnr9ELh/G/47/C69q4iCif4hDcWNPYSqV7ghT5DshEvK7b+2eZDryC
Z5bIaggIiLkUYC7QeQLVhlfRVEySnJQC0D24P+lD62kWUWHN2NIVQbmWOAqfbJ6D
JFJF/eEpZnfGIrWmbsrPgarDc4Zc3fZeUiNxXAiTBzTO65mNSWFpFDvztV36O14Y
Cqu/bMK+sYaRyLcb8nkEtq7yAE8uIvMNqIGfr0SWAS9iidKa7wK9CoPhaHBqNYI7
zzbWadstmaYd3WDuqp5V0sbYH+7nM8T59CZutP085EB95ileDjKXjlDo6jplsA41
N135cmsofuDI9gLEGkTxtjt5iHJJPEo9nqa/LXCVO5oxJ4biKkCmXJN7P6my+JAh
8cPXjwQD+y3W3NNY+jW35iy8RvkMv70HYvhpkMGhiCZF8wQ+5nQBEnt1RPvHzZxf
t+dU+HNjnOwWq9rrKPR7dIInXdQVVoXIDqauJEX0W6TUwSwgSFCkF6UHnFtTjAPv
dYthHOZhyh7XwoT5F36ByAp7d+2Yw9QG427LkUH87LeSiKCsmoE+z7uU3Or046Lx
lFUg7U67ANjk+LRWMtrDzy9j/1IV2at/L2o8udDd7xaV1nTv9BLIKYh3yywjVJ+x
DfQBf+apTiNVNR+w10hSqyC2y7vCAUSa8ST+xPZJPY47Std8Ws3yBLZlN7J9Cx8k
4/+vagP9bOqDn/BGPS+N421oc8y6dMBcpN/IR5XEdZyGf1vDRbFkLvOQEOYiRKiY
Ty0VL/aMVHvOcYCMNoSaDX95hSUnmWiJu5Jf0zZEQnXuiwFQltLmcEOGSn7p1Av0
LwiwV7F3tP6l98FIHbmTxSot8Cf6cVlUzbM6PrY6Tg/S3j+Y0trYIxY45nYmgMiT
o7KnrC9AHoYY8OlsZoazY6t06apgsDsxNF+xZjx7k53lybE6+I7P89LVjrFnumbo
5jRdaz7W4AVbeqkSGVaj7kf1oUdihDBmiOSijuWPNPh4a5iu3/LKQwYqr6u9lFYF
Zmu2dhnNkz0Izy9PBt+YIeOAu/6QxbC/vhRmnLS7uOmPebEV5P3CZ2yVIgs4jv0k
Coy6pxi3YY2AXQs6SRtxbiO9a9cPRoADsSuKTbX9Ds1w4hEuotnP1dcx202/6xb8
R/MrRJYfOOd9vrpYyJ1sy3tFw5ntl25B6JAYnErnOsE+YzQjDnPlCFRYkJeXFsa4
XeiPUB4gdby+bhHdrC+Jo17hYh6aWrkLVckR9w+qX16CVjqWzwvTy+AbuI8C339/
FRgm2ZGg6VF54tcQdq4xg6RRh/YZoWOoJ093q97+SKTXg9HJL6BXfE0m0KfmEeCB
KvQSYOYQN2IwRnVpyIaue84fbLckTpNaEYu9fQMrs4SFs2cu5gtdevNFx60N55ht
RIgjyfLJH0XF8kP44/2YA2akWUmNrIZdG4r4E/BiG7C7v9i5Wro4zNJPmpQUDuu7
EXrbhLa9UhxY3H9dAYWdmIWkQc7GGEWam9gMwUtq2X9PHDIlFBIMtA8ns8W/uch6
xqiiKxi/kDlJW6e1FkoXIp5DXnuS9XkEcbxNS9aqvQC9TNFdGxDweaZ2bQ+rOXrX
ag4yBSHyg+wfDIa3k3qD5cZpIlMVe6h/SD9pJwbkUKmQIhUBYIgulokkL1+OFVDR
kf7F2RgfE0+zw3TFJ8194jCPQLLCl3jT8LUJxX3TEBDeh1L5v3LNNF33hv1+bM6n
ECNPrLKlUK6aqAuAr1PcyfWIW2Kesuej1ZNJZeokPEdbLNienL9IiToMEk/qWjlK
FDjBB4pVfFTj5kSpVJXHm46ESPSEnXzbb/8tDHlj0tKqmYoaGgyhzE5JGeh3nr0O
Sf0t1ftSCG6XQn/cMqnCZr2VYiqlVjCbcOiK30e4MYw8cebPgj/V5DhYKjoumrJr
Tq2AK7ZpHKnM23UVfhMtwNaZY83f+xxvZ23Rfo3M02Y6eQiymMG3I+7n5Xg99pxj
64h/h0brtp2DalJOxgBsn/lrOyVYhI8OwzaZRQTvM2DXI6eNTQ3ET6m/H8ivgLVl
Qi4DzPj4xK8CC4nqcZnNJc485t+F7uH3aBehmxj5CgT7ag3l3J9NEBLfd/DPeAk+
cr1o28g3dJEIMq64Y122fDZ4EeUd2T8chxWUwqvoofvIAiJStfN6yuSL+NUB1a0i
35YdiEB1I3j/ntJU+HOCDH+IJgXp3qzXOzhn5q/iRX/yt2/XAqrJ4QEJaeOmMEA5
2P+0a9MGzidLGwHxHYzdTHbc+BjIp7344IgOWSkvn4cRDCk8ZlfEPY9uYE0GFArD
QtQxKfog9i7nMHPQwWebtOm579BCnneZi992Xcy4zl6aLBuG1BKAolv/nqD6PXfW
1TesZVN3f8Tn3BkIh/G9cLV5mepy0xJpxhq1h8OUkXPic2RSOrXaoqRITsTjkpLC
4QZUeWcDjm8pDKODxF8lZluc+VKYWBIjKXkmlgeCpMWq1/cLBUZpeGK7sX+9po7w
S25kYp0nl4w6yXZpPEWbf6CJ1ackS/V5Xnr9Jc/PeGy308MXV5/EnS4rx3dTEuy6
jiyjQ84y4JGXn8BDHQYR/6Dl9GCyPQMrnGYugFRlvfROxuqbl0BHt2W83BGkvHDA
eGJ7FpvYVTPIwjA2UrbKXU88xTRY0KPW5Q/RytqpXPXuIktDSouoaxV6dnnOC9vy
hilfaO+0AK6yRqib8EE0k1YbCSG4mTwv1Gm9LakyHYShhdjgJDJhP6Jtr1UQHcqf
7fW07OZPvz5EC8kzxYIk9iX7C6CkpTfN8fQYURfDb+0VogdDV//0iRg37wQdDlcW
zYIOp32wTu3iMYFvMXEGMu0LgzwL/KubyNJ7qIBMyY83qkQvYoksg4w2Xn0UXg4f
HaoqyT+Cfpf7f1ZCEtwwaQY/+9b44uXSZtVGXUfnRae6spgQHTMGFlf11bRsuQR6
UHhvz/ltwuwbisNIvZ9jBKYmu3Xj52y6NuzWCmwvTEDs8HZEeQ8kcfl68lz9cc8H
glSqoeFLeZu+hIy8Y/bLrJBa5v+GY7/+0rUkonHStjqgcrjZ/owQos6Tb7jBg4QN
drlQtxo5I2VkvgBtAfOHXMfvggg2f28+EDAoO6aiZ+dbLYBnlqLIgaLTwFiE68NL
pHz6I4iNIqqR6xVIe8cAVlWo91ND5JRoczEv+81RMoPZe1eNW6UV/xZHKctNnLut
wbLOkJpGJijt09WTEp0KhzIuF7Z9NV3A3o0RDfSG1fofArYCqX6XExSn8rJ+glzl
tf/PUW73hATvLvirxYv1H5txLdzf8flRNIOb2zUqpKx4ihzUAePSn2ALfGH1IWOB
BJATNhnRD67jJNFtTM/d1ny2IdY1ze/evTljttMwpVZlXRduZRjeU6s4KRezh5oQ
fsBP1yXbt8NUqchYXDquuOKusnKTaWVGQv9ThOyUvLkKtc7lnZ5zVYYN7Lr6a3lf
jZgQ7WJdJ/Q6/ioY9tJeRU6ElnrdUnUBB7qHKxZkiuqEoHUiIjJh0oE6nHlyFu0J
vVwNGSLOOc+afz9r0cdUuWI+WZu/fdTOL3TQzr1fvCGGTV3pcntjfNhdlheTeJPP
3HIH5Qjt4SVlM+/rhB5REYApD20YH/rXtunwwkNLcTJWf9EEUyH0jR1WbWdcy0vy
AHPwAj2ISL8o0A3iAiZUkWQYeKb1tyUt4BsYBM/h3+ycwNqoAeOcO0/QblxMDzBc
eQr9fzeO5a8LwF5ger8oAPsnc6l3R2Hk1uZMDCUlyUpNV4p+HP92z+iEFf1TVsIx
FW8V4jim+f9oLtOojjVe0eIdkuRH8AmxwSJpQDWmtzPkn3C8VPi1QvszZSmA0lVI
Xp3EBSPBP4CJGHq2fWTcQZHKeZI5rIwnPVTH2ELHlbcq7+v1fETbQNLUzbv6AuJH
TR8thL5RvN/Mofl0ldMs9WFWYaySulr5hFbvSp9U7hhVQyM7AKA8WAPMZL+WQfGj
i8ANHVa0e3C+KNJGWyhU1fRni7kwBpzzrRlW1qOjVUmJ71O4b8SLgdOfrPi7El9w
9ZiGlAaGGfcxDS3K5e8vXJPltOjtmO833d+dpJnwQ+PKSuIu/eISvhJCQImr8xoc
9nGAToDbXqSpeDaMtPur6d3/Hh5h0LMsaI4yGb22Bnq0bguupV73/aSSA0JN5kTf
n1xmyvBIyxIPFJtOFabN4XZUjC/yfXxxcxiTuUi6iHmqPgBqqsgDzevM6PXKKCSJ
wnH9hsDUV2v9yhD/qsRWs5xLp2F13IoVrAoGztHNMGeaxQTpEeeFR+fH2tr+sqr0
JLSesjBDhsv13uBSaTpqjMVf53ONB3KcWXnbaeAXmgH8eE1VpYathwhnraMLKVi7
jsb08lwKcTtxJ7KQ4Df9T1sq81Bj7Xko/N+SVAdpcEFCL2VR2fTCr6c9RBexhgzd
neiBJ1b7Y8mBJNlllaE51rjo1S8cbv+WOEJ/ptITcWQRfBuu1EY61ukiZVM3CkIA
G9cFIoaP0GQuEWmloHkXUrkDCXQ5BK9rtulu/rpc+bjX/oycORxG9mqu/UgIboGF
i4lxRL5RZf7FsJHi1cI+UttdaCE0+cCIkmeg44vy8HRgKb0sS36Eu7vc6xfz5sK5
7LbzGvOKcP0Dj4Lm5xCnsScEH3eWuRDIIFWswH1qrTgioLU7Wx9Jf5JTNFfCXqcZ
3zYUycjSMsdoPD5LB7LWmCIz/OtwhUWRePbRCyXztu6uGhawQnVLTqr5lvX4VUnh
4DWSbRjX/qCAwyX41fZtlYtnPjCxfWz2nxjhWBJd+CtrBOxmt7yTakAQPo0eQ3Qr
IQcmuB/1qoOtdwiW98VBY7pGjL3B0RmPEcwD43XcyYiddLUO8v3k5SuBRhRiXeNb
9cVGvHmPkeIZz6OxuszaUx2fMamcy12RWTk+4EBvyB8bOhUVrR0cFLvZW4i5x97y
ehF8fkmZD+HeHaBenWvl2mOygIEfRcIh9Mr9INQATc7LP2cnB8XqFrEdMtx3CoTI
jgnqiZy+YKVhz6V0U55RY2Bqt8OVsMGha1YDtE4/4os8D0zTQEA7KTjroCtC88gh
zelpxeFEsgUswT0V/FsDketiNZ9Q061TC7TKeqzSN4oRE9deSSKVlw81fVpKfmi6
jUB8VhCmvcvWMDqavg/3c0IM7o/AJx7d+RwOYPFrIuBwzF7ZJDk6XItFMTQ4l6lV
OljqU4xH7gxxOa2fq8zy6U01YZY9HGjFq8Dka/t/VOJzacCc2x/g8o34jimedTAZ
vWtDhSBsw/06YYx6Pnf6p42wqDQ+SPHPyr6gLX3GPxqfQ9Xiz4vtcXeDAqka2m8p
GCdReHZA5ZTGNuYUZYDU0QQ7e0np+NVg58V6wK5PYjMUx80A6/6ggXSZ7clu2rQC
mVLSMdstTOtM3xtzNBAjKgrJ80+i9x7B2R4qnNYlFrP+OXaG4pCviwj0H9lyJFql
LBj1ko7MFkVy5BIFK7NLZGAJGfMOOLEKRs+3suE4wBvPsS+jkIESGv+PySIniK/T
bHj+F8f86NIPvEYB51HTiMCPzNsCnA3aihQRG+T7TT5opZtlZiT6dB0UIpcMQvAA
53wuHqURhA1qWGEebJp57fjKjO3sdREEicgrQKk86Gh2+0t7iSRZk0dbLr+XDykP
kFudXtBA8eAgmX4RpAxfkfE+QyUudxnKFYpDrPtSuGGmDlkUdYhydrLLnRSvjniz
ba85rjn/QdjYvUjamHmzvZOi4+NkowQq76D8huYhW1XPeQuVQL5ZzyBnZGh6ilix
5IdAX3oyQ3ntxIPmuD8xwaxAruqVqSRjLplqP4LDrHMbVsh/z6dDX/+6NJtrUXn3
CKIm2hhin78DN7WAELPYyaIi9s3NrdjcT1joOQYrFANnI2Uyka2d0RDAE4IEn5/W
XszHcTueNAVZ6La0U2nr358/8lWIeBVP0Q+2jEWDPo2fKrrsSY+aWRz0fmLzdUww
XOfRqNBMSa+n6vZ/7JFFjoXm2mudiq02OQWFv8hWAQ3YuoCxjohhDkAjR3SmILTA
tmm26HC4fJLSKUhqW2WUKE6LvF+i9sqaWbWuEYndScQcU4R3a/4E97le5bMNV608
mQzlN5UruFHeAmBe8aWzwg==
`protect end_protected
