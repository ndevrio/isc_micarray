// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
EV06Fx09uRBHvETU2J7xmwE5Q+Pi17Wd84n/mnRt9MpSuuJC/VdFZCPhVkBE94Ku
9xProhCn2UeFxqYjba0zgr/bQp5kJhATdyNkjXWnQc3UT0171rGNEYy9V81ydPZw
eGmiG4OaPlUmxd1wPfe4BE88ENrZBPsdrlPX7ObVd+gQ28JQ+g/paw==
//pragma protect end_key_block
//pragma protect digest_block
eYRy8N0s4JtXXjS+fIqYjAAoeKw=
//pragma protect end_digest_block
//pragma protect data_block
9WKehnTS+PyP3MKk5mQBJ+5q6qv+IZ12Z/I0UxYhkQpSCfDpAXPNH6YsHb5ojpYQ
+a3KQwC8Xjeol5yx/iWuWJuBfRL0LmpMsfNozFDumeSTJeH13wsphbGzC2XONeyb
RqfjGnK1fcmUQpV0r28occUOLjVj0yNdJBwqGLTlcTKZ9xP6FHIoi+xKBOPPri3w
hM1nXyFdbD52fhwZGJsq/AzhMSkX8EC05c8Fnn+1gbUrOq3oDwQno6avS9WQL3AT
ZDH+z3ET3Vur/ehuWb3dmPunJjsrUf+2YfDlm3PRUs2FJG41M5i4X0zQ6VwWH5a7
EW6Z014ezgT+sG77/JC1gEi29vzULTb3z3ewdyx619x7fXBCkWCeYiBplJe+AahV
TXI8vWdZOsEE9rRmchc86QgsgW9FULzvA4VkAcAdxj/LSetxYR8Fk/u/4U4igs/3
ZuZzALxATHVtBFL3nMUPx9Jw2cKyDS0bXXeLSI15nrTvDB+OCiVP9/o45yRps814
SQwdRxRw+/OEOhc8Tgn/12ROSWPTdqs/42PkTNf7s/3IsMtFph0qPWn4ikNChMkY
36chEvSo6RizfSrY4f5piB3LmY2tysJI1tRaCN7Na4EKNhL2RelWupLtYmInGupM
zo4gRlE31Ah6MQTNb3kIcKmYecUcCfYy4bKLE5olO0LNV5ITF6d5LHfx3AjJZ302
IxjvgHVreJDyu6O5Q52Csc6/VX61jz4nAhGcKDkFSOOqHHIvLttdb7QQQ//1jTAL
6UjC2iRdTYFke1AALkwFmwQghX7pQnz0vbziAy4tR79bgQVJH8eIFd3YwFDBgT5g
+c0PGqTANz8cr8AkyR5AcP0v7S5feAd5oo2d5hGf3lDfMh+DYmjYIHEKWfHqRoOn
PCVJwXr+sNkP+4QiWZ3mEgAeGrsJgKOu/Q2ZT/0CGGSVcAJqPb15OOew5J0/aBWO
tfbT1/AQQ1QlD0bJobhhhFteGGQyUw9OFJSjEcnAMSdYwmNTSeaZwwzZ8ORIaiZu
f0lktILQtiHb82N10hI+XdGGLmaLGy2DSBLItrRUJl9RbU/AenyN0iH+7dDUEyem
+D0UIijRNZO1S4cmTDu415/FAmmDzjwbndH4vHHAA9XtiWzYae+Rj2McfC+9th8N
1FJlcGIJvCXscPBCFr9PB/fu3W6L3jVTTB1nI7n+CC1Gkru30p/8t8CxH0X6+29v
7LMPdcNwyhFxXchcRp+ZU2u2xopJVE5pKuD9bpDSrlnKMmALR6iteJtjdCPuySxJ
K5kIga0ihs0oomGKEjIKw0ocSpr0Z8JoD5Sa4PUnQQbE59GBg+y4N/kdiP54sY1i
BAHS19x6QGWiET7Fa57OplaaLanuJVgiFC5X3bHQ1zV97oUTw+qa8ksuM3l0dKL8
DbvrRb7BaxgI+q0zliOj517HKCnZp76USO5OeUe2t6ICFw7PMCZY9RFXuabNsLrs
mdNxGC8BZncc+VFNAd3zrbeUT7tFJirxVswTCpfnhF8BXlHzBFKTKtoqu76IuidH
jQl0xYQ19nEUy7OLecyHKwJ85FXEFbTGDYa7egS/hyyBSgIibrR6UUIHsbAbbIGn
0Ln6Jss4z6zqtjfCjZB73rBmGFR5aUrHkpOg2Aw28CO/PhjB3ek82hayFhGo5CAQ
/Xmq0D5xVbLig/syF967K3ogf5BAbxAg/Ixwy29znSuDjyEBDxQbOR+JaehpJ3yo
jVOiKvzrgqgNbX2VCjI0by135Yf45ZddMm1wVOT9v7h5lQhVxtFSLe+U/5PBVgnj
eRjAZKYR/X+vKGyNNbIYS0JcQxrYrPojNC379B/izGTahZSLCoaGVHXD7rV/LM2+
JFlAuMlQdhwK6V+ASmVbHhcj4hSKL3MAtLZk5Z5DMR39mjokiGAXJG4C1if8A59G
rzI/UN20vmXVhZQ0ZPlAObk2AOlny6MuKvwA8UiYROtXmB9HFghrDh1UB37h8T32
1WACS/HVcg9CDaaGmJzjsAjJ2DZzZb31XFGidEmmku87GinM+qP17zOaNdYKuR/8
3k5/ZiUkUFA20/jtypneuCaeTVMIl9eSyoXfYSTOgeaTIYNLnVk3x+wm3pQ/ogG2
o4q+1cizTh/kT0DGff1gK5IJNQ+4O7VuPOeCfsMiMQWHMBtUV50LbOMFR3hkIgf4
zCkbysPyzOr8b1+IKa8TFMxbkW+XGWc213w/8/2ErfK04dbJCXILGmAS+KjsEW7n
1JEYp2Xab76ullOipRau56qnroF0+N1XaTRNR5VXo7CxtiHxWgfE4nc0x0YtW8Nb
E2pDZVSBSmA6NI07Vo4Rc36L8MpbGzfl/Qipp9XPvajXRMDOr/YqBZQn59qxMhZz
Tus80801W3ROI/lmEZda6prYbScQ6VUMCOG7TIJbEYF1dbgW3xrAn3NEf/dUf6WX
+9B76XPJP8pmu38QFFdFLQ35ymZ3Oa6h+lD/gPxbk7LELcujyB0oyPzU4lPzl+YM
lPkPO4IxuBz1or73rTrm2oFTd8fxrtPNTen9HhqlgAMEnLBsayZdyZvylNB2l5z4
7+epy62vMF7uvYvVcU3pQ2uBYsEzEmBuRvl6j8AVqrMR4x0EgiUijRusYa/0b96o
5bclH/QXG/4OiswJD6Zve6V+RQIqMwOcd4KztRQzMQ8XOcAesXXzxbEOR/lWe5O8
HtHc6w3YxF0LQouQ0bTLKDcB57Y5ymDf85AmpfE4OG20xxd/KJZYQTDCg4vCC9yM
y9tTnMUs5GpwCJtV6CsibUPZXDF3+rWklGJbr+YImWtvzXCEXygKz/RNOJXL5gg3
8rY/ywNcbNqbZLJ5A39XOZ3Kqm3cPt0dK63UufBHP6GuOcY0smKSAbNDjMOoKbhx
BFsu+eHdGSHq0w3OGxhW+I+ZCqhqC18eXCd0hVH53uMP/rI/Lkr3AUF2PDHmkBXZ
f9zGSIqqr6JpW4gZlzKfetBkYTvsB4phP5tZyh3Wl2cHOWLUG7yLkK71Rk7Z3p80
u7zm0iuQ+vKbdxUbcT1PwNvs9F1s4dO57t7u/gyA036BpnCLk6aer1LVDL/lgibh
t4OVU5p6QH5VytfuBOO0E+XYnnEXpUJtRbXaFFpLHFxd3jXJmz9HWW0NgoldcmhW
LKWgm9dpUGf5JeHzdqqHPa3MyWhiVQ/vSOU0tXD8dUdOK576bmURG1Fms0WqPg7e
9z6tIN+s+PTBVNPzauKUfMmA9UZnNtH1THkt6DNNRczCHx9YEzoolLAEVrB1bTEr
VTm9oSVheguu/3yrgGGK2hxPwrDWtEW2kMbCWyb33E2P0Nd5mqVfXEJ80MZ/0GMV
xFaPKtGBuSvFvXT36c1fW9/eG1VPQROk0TUIi83g7GZyPOEUVCbfCrns1ykyKsgC
E2SsRHyF9v/qeExuJMk4/p49BkbFQx1I8ystOV5u80E/TkH9FQwuT/NQRQXNXcVC
23VGwJZrjoZSBVbAcmv1t/iKeCmH/B8C7ITV5F6Cm92LAqMbXx97QRz5TYw5hC2j
3Uhrz8mqzLkMqcbCipADOVr7nXbuidRFRiQry9oERKXLfMdVWYyQZnRHAUaojEbM
4RbROcU8UQVZyzWCql9dL0hJNf5t3yJRYkFqTxTyAf5vKsV8rCu2pGHsk/eTtw0Y
n+SNn+100GGNG7GhyAmBxppOK9kmRcQ8jxZcgNTjrbRhFp4TGoJh8c+g26EKrEPt
7Z3Oqi8Iia8c2w1jkLQlUCxDV+XAPsK2W9t/1GO5/Fr9ozk2wSMjrZftJQmMMrwn
Rb1b3sWwuUsHTML/WfbN3f0Z5OwggsdGeBXFACNB/bjlW0a9UXgYCCPgb9CLM0xP
jvSSbLXiHzVJ17xYx7D/9d4olWrXSoWOG3MWsMaZlVvLruW/PghpiK2P/XDWZaOF
BE4XTYh+iQrYJbkQHOPCHCivYu0MZvm6UUOlgMaOP0hVLKD71L66Cow882A/S2PD
ZHVsQYXxrrNbZJBQoNuphS/IogHeoNcrlmkW8vS51YHYoOjvFaeWmbeLpvW/fQSv
aBJ1AWNBP2oDKk/9XfcvNIt2ocpYL8IifRmlRWx46nAh8au/SRbtVAExhQUrNxY9
dFlVCRDbuCXn+9Y/aXGWJmkjYgJl7W9SuKH0/o48y7BEr4+kaE13CWMaSy8nnIx+
7p0ei1/pAUyHbsOj0R6+AUXcuPhbEvy5GE205Cuf6v7NxwLNyRVXBVH7X06FZfK6
fbyV1rCIL4teX+ogEeaR0LYAz9uRE3Cn1E2WpGHv5bHSUZcodZpKckKHAaiIgyCy
C+fXHQ34IH4+1/GZplo/fdYITwCmW3aKCe8Qq+H/BwTKWy73E0zwGDZlO6p7NHjV
/eRUShJzRJS56FGu+hmU0OSfIYuxIQiCKnxPjTlV4TBMikjk3w+UOZ0SxA+ZQ+3O
bEeWu7nUfmd/pQeA+WxfNBnjF8hogmjNTfDRpgVgNL22OltOIxWW5RODlKtyhXOx
SUnjpuEcOiFQzzZwRVy9ItqaJsluQZKpvbaaAHPBNOAZsAFOpCHhNmefqoTxh5gB
0mJEwPmnaVag0ArwI8rhFEXE2vC1YNPl67EjuBeneRzFtey8wBkl5hAYCDdDYC7V
hLVqqU2WDBbNKkncKRcP1W9xB1/sIKqjxyp6YACWvjkdLCPT9Xj02v3tovPSiyPu
6FX2aaBoGtZI7gHKFcusNRXDgb1Z2n00xSbU0Yed5Nx5dh1idgeI8jeK1ovrTO0v
DF2M0WBqQzfnBkLaW9QhBBSoxClmAnPuV6bxxoLhQ2X1fwc1dneME9dFTxBsvCWM
efrMLmbtxzwWd9G+BH4/4nBYB++tBGCgLOMwqRAnMGT27F22ac/CV+8LjdbZs2u2
tR0pupJuO/ogTYjLoAbAAaVQBm2EYsdK1dgs37kqz0nz0DJAcj33AgvnhBkgWUOv
/M1NaF0gpJYUrDHi7/atJwa1UmXEJPS2j88z8XI/DjEUNFiXpgsNpTiGCKPvX6yE
uO8SHEgOc5UvIKDVt4OztH0q8kK78mM36nItp3MIxpgjcVJwQR5nKtiuxaA6uxUX
d59UZ+UmcZWyNmDZX4gq25mAGkzKxflD/32/20EcacgzzZ0plFN8RLrWn8SwQo/O
eVoAFOJTVglHeHAVmEKfIBxa3LGIqHFQC1glcSlfVP5wjlyoAigAh3eUnXUUoyQo
t3jbaU1uVwH690YdpgvxFhEkqNtsWZ4vsZfeBPyQfawD8AaAqP3PJWT6VcCFlHfJ
f+FKY9+ETnQ4dWqQz3rhZx5fqO9CJaY0nDWaYyCBuOlJQEEfn8hWQ6LWTnS62obT
Rlm7ZXYaSRPTM/oUZScomzf6vd6M7scPgJCSuZkxWvFlRS9xbC0rybK56/krdxCz
la84jsjwiadkmNPUsecm6zSayfss17tirZ5wap6hexj/AQI4m4yqQslAbhf4nbwf
uwfigjIYPnIZ6L4OLoWDjlezJdkrfod2EjQdnNhAO0ViWy7WHHIRAbhdkDDPIvlu
h55Yq8lJhHa+GUp2P1zS2Z1I6IDd4e6kzZaJG/UwRTgjPH23IEMAaKid4w/FmzWE
EoNARxVxlQzJcEV85XiE1eSUvUkt6ZiDGChuVnd7m/buTjpKCOZMo2f8I1zrCsim
13ZRAzZFaMcr3pz9s2PmPp+X8JXPJVxRvDTHZ3N7dJ2hfvhjWGRbOlDVQfGTvvFA
hVkgZ4vQzY7FSlaq6/zGQ3oWfIvb4oIya3lDSolLN/rvZbGG0zs7atIoGTgUmoRD
k1ESWfcwan+RFZ4+Ow7ORdnj/7KPvZUFm+aU1qJWxoxxbKV8Ws/PSAP9xMz7z0Rt
lEzUv3RpxkpcKSnJuzwmPKxp5IeewfbCfJCoCN6QijEBBkbAQ05g0Zv7r95R6f5W
urWTKr5wa3nMoDUI+6onymRDs2Z1J65gjltQf6ZvR2daLPS+dvh35evk/ggDg+AK
JRaxN9NneJaRFTmDDfYVOgrlKXgfw7YkC/EFmCVEsGXJB8d0GiVfjnPnNmGva5YM
AUzIW8g/BIKUu6YiEftWGUNzQPhA3O1nyMSP45rJL01sFleT9npwk+b+aFWjJ2Nw
eUenZ03gRLF+kmIWKBRgshxNDU5l0Vng97sUz0WPXUuOT9ZC0dHyYyNTyW8as7aR
DQs0XTpay8vchV2S/030KM4hNigtk+Z8WhlK8VkN2yThtn1dSAKAQ0Hwa1Ub7vQ/
L1qCIrc4yO1QVv+OehUptX7f6MlRmy3VABX8FJ4N1beXoLrZLIoL5woPhCbk3cF5
HoN1DTnLSYqn75Dt5nugh36f93dAOhBsBPgbMRsKX48iChR8Q9nnxjcniTNzgJ46
KO5D5CMsumErqUIOdG0xQI+OF01/C8apo+JXbwHED0UjBmjdMtD9cK1iSAXI2nrm
/Cv0qkXI3LkmILCJgK4NDkFKq6HQ5n2o/vbK3YJaAbEqwbbImiU7mAVt7TZCvJnI
CEdkD8VLr4uRWP96R2nvT8nfrPPRBuRzrnK5vlsRgqUUQkbQG9JN4rLR9bOLwuHK
gMACh0E7zUsZIBZ0taK9SolUxhZaQb/73sz4tmhIi14MWT33hnzLPjj/t169m1uo
apOP+o2TN7NhbuAys/LQmRUu4PrByb5NyzuY0VTHQNB8yjaLNSpiQQQyxOj3Jp2B
fLwc7wnoCJGEyXxJ81kuoNgIz8XZxdQDbyCA3IteOJGKDIxVsrA1YQPIoH7zh2S5
EJi0022LJZCrcj/bWkGIo+H9Of+SYWY+vmktzTAeVcbCGhKzAyDmuXvGdXYzMISB
D0+GUHaiEaBNuhYHgOLc4fDfOdQoLGv0/2VKO6F5zlwp9OAo5mCkQsNBwCKEau21
F+Qf6QCLdkD1NX00T2foj69Lx6QQqvy9PL/QKl75HgGrmfMuhLzapFUGEz372cjB
HEwLlV39f4cVizsn0Dxnuzg6BpGBhgtRMmyy9/d0SePutzMfVt3P9wAX0Dgn7uR4
ttoZN64qQRTvyGvzN6hpaMNGEbfOFjVlsVATTzJgFrkjARt3ZRHsxixfC/+/kOwD
9C7mdGDKEfaYxb6lkNHuTq1wbqMQpIEmJKJjiVCU84/iNl049K68SxFaUHRUvOuj
f1KwZ+HiprXT/4Tu/jaN57Fb+wBreDOnRVOi1kvou0usw5FjsGpfGoMKu5oURkxg
9CJjaVMWgchVzZrHjFZSDV3NM/ueILDxc3rfwM3JlSFwp8RBy2tP0qKbNDdFUsFl
hpuwpsIXXJQSFkYWiF4AL8CAjo0Sy8Lo021kIlfQztoUwNkF+qgZWsCchhH1Hita
Q4MHmzfYvG8icB4xv3WtKG4DMJsNq2Q3rP/5zfAhwwcrctabRg8z+Hm5kKj/MHDI
jsPZZE5HLFOaCCRvo4vVKBGpwWJoRzMQTgE5gVsncaWhmg+vrwPWj77X1YAdlOAS
yCeKvLR1VIz3wqFI1gSCPLlUwMerGuLpTxqckQ3FfzcgfV8hODtusTCGrw/KaBmO
CedBkOPca/BsgFvW5yBjsIqW3m6jkFfJp8IIxz6G07xakmHh+cIqfU+3r+lFWUuY
bpJXmTFRlwHNJUzWmS5RMKyBZk9+y0uPlcdkNaGFE4QzPqQsEKUoBKbSKQHxFCYV
Tfdxi6x8XJdWChEYI4DnBOG9SvEv7+WEXx47MOiDosEOVC5Xat4ZA1nnyGlXsRkL
MPDkZYK8+rEUswvepK7hRlcQ5y93HKm00lRDJ851arjnAb0pgQK9u25QmCl/eOnN
UjAQBRJAVGLZWra3+9bK6OeXBqiQ3Li4aDPiXDbadAzdPcsUE55sKGnan42ud0vc
8rHrwI7Cvdukwn3EZsjt+9iVRJEur5LaaCwrWEGefALcYacn9hQEsfs3VZXmZvxS
0lG0txmAqypn2o/8szXCuDqVd5bHSsTXF9J1HczqbpaU1r1AvB0J2wQ/LSH/3OMi
cHvO10X+4RedDi12jb6ZWAzhYu+QcpWuelT40oo4HhqB+XjsSFJZrhaYgqB/0n7A
xqrQrMo1VJGKSHj3oRp+0ta4z2Oh2f/2C5cuotILyw2J/vNC+F2QM0urz5nEnNW6
b/3HxnnZgCpA64ym+DrJY3NzPi6gHV/X0VTMKXPKy+MC4LdS6CjP3mNarD2TnHLp
m9e2seTFBR8SQQNPy4TegcFdrTxTm+VoHAsLGDzv7LzV8cLg3IzQSYu6B++g7wzt
PwGlHVdx5QTAd8jufJyokMaUxAIXWUE9GiSrkfy0RAPpi8DOBK8GBAFcD0EMlOcb
WCyfiuGy9F9BOn8itNd1HGGZ+o4X7s30T6qGOi+PxFq8JE8wt7SMBwwl2/lr9dyg
+QZCLyi95Ii9MG1oWcRN44kp32epx/RgBMw5MyBhs9F/Z39uCAUz1UVIVOObwa5j
i6AeSevr/qNlCMSomMUM//L4wF4Q6C+sJ1IRwd1mUpqTOvCb4nC3CTvYReEw4CRz
z7TtOYQKDRUze2Ugehr4iJ65l14bZTUFQGow1HUwkWMa6kokm+1+BrH/J7tsCR2I
JAyypKiFQz/HwBJQhIRNq5zWV15n/2qVkWYnd+6hqu3WgAAa1egTvtZM5NFZTZ8Q
aWPPZ7/9x8kTBMIVEAlVKZSZkdJZt64ozCNeE1NvwewGmU8Xway/RvNpHAGxHeGz
AflMIOYitImjCoLVx9Grsl5EdlEbY6N+z0rwwwhNEvjrU7tbXLaseyiyfuZe17Bv
zVjCJr1KmrV81p+krFMy9jAua5Sqrc3SJMq5Sf1XLYnyyJ9OLw9xYznvSNj3IDth
PsY0tSuzJklWkSBJWedSndTPilVEUCoHat+Q0aE+U5ctmMpKQNsPWs4PjojW4mb3
m1MJ2keqqwJizqXuvATxzjYjtoK9HV/fGZ5ePipI/LzqoaL5R6b7jNvHa9MxWZrv
HrI/39ot9+0e+AMocjayDhaNq0W4th+q3zxU4NmTMJg6pBxOI2UiMkMRJZ6/k7uX
/9nRIsVMpAI835uggnbmYGxeJOaSpqH9ndc03eVycYBW010tggswD4uZG6t1RlzC
OH6VLBEu8bUfgRy3pkB80cdIR77LD+yDGm1amsWSqUjz9IJRoEZX8s9vsWWsD7+F
eRepn5PUjeuLAJ/JIIKL/Z0GCpMDqJ3fmm1piVPJN0fiW0GqRIHnL9fDzRsANzT3
45BQELXJzVjLHs1XPgIlVN2qj0/XQuZx65I4si9qxZH1N4oP+0XFVV7R5y294rWn
Wf3+58kqoIpg91RSab9fSBohAxoVGoxMa7YTbLbapbYjylCSkb+FSe0zBvYJDVNC
Ov4D7X0FJ1mh/DUQRioD7Dii1z63a6MkPLimXXoGUAdY/DBl0QBJZGoydtbS9r5c
l+q4Yhs/kSeLyYummetRW4tmEjvtIwUGBxD3KOv2y4cGkRYiSco+b0lifGllE2l2
oT8mIMkwQod0neBlo6bOri+94Mfu9IetOKwgk/3JhjdeLqcFrU/zvSt4ui9zMpzn
sQKMIGdQZP7d8/SFB4bUP1zALRe6YkODYuILnIE2HZEcThPrAD/jTDFDTZ8GqYKn
3FaQNvnpVebaBG7p4T4ZdwtkzBg5vqHq7zoJTZj7X31UGseJNnHgSkHh8U68yagj
Bz7UrVTYP06vt+Ff1tjL3YKzgltuqdx/eBMTBH0dUBy8tZ0adroOQvF1rJd3GBJk
dMA0IDfZTsGKhm5m2noCnD/RVatrCHp5TRVTg4wrLoEQ5RhlKNtpRX3j0iy9lo4z
1NaCSQf2mBeRK7VSE1F9me18HpI6n8ZUCXGPefio/b3eqUYskFQc0JH/VBJ/PZm7
M7Ey1h5LNbCiABAUA88KyzXoW3kHW168daWXUqH+gm3l2e0aw0dYfWinhoM8N22o
ctQ7AGbi9m6kWb6JAINVLqUzXRjfVct3qgTFPPEIgfANb7BeJW2kbZUgV4eZmE4z
8yxs6aYEbGBB+j8Zw/ko5eXWOOgBx+OQ5DdhIrZEeK8iLSBSLgie1jaR9DITTuj2
OHkNfR+7DgPG2OFJyWWK5MU1lcQHy8fnSev1kcqQwJ8gcI/jZ8ncR05gkvEupKr2
RhY93bFvD60YWMO4v05CG1QGQ+qOEsiCobx8ajrsFxilSdiNTnu1fxeRo/ZC1O78
RLuYpNTu/i8984CQQnI9mKR9KW1/WZmn6CACZJr7cE4UfNi4CJHM/nbeCYsuI/Vd
EhnFOEV9o3gB0HGImxcDbKn/ueaOMSXNtqPnjE/mMaWW6iCkEMV08pnkRb7zFzMq
e3yMmjoOfpZL8hMPMvMshKkhkaBSHfQET1npatoR14GcdNCQ/RXI1HxTyy8TkokL
K1hHrJLzsLIyzYgaxlaxTtjEdySu72Rp95KUcWvqkfS0EbzbUb4SWSfJdqoES2DR
W0+wseJanxNSTIyddazf7SmN8/tq8M2XRMAaf0hlzNLhodc6jo4BYrosCpq23yXl
4ymqU7Qm+KxRcgG/Etr857ki2ZVEPHSdMYQNZDqZvjGi06+bDTEcs0sdnjZdrsga
6Ir606KnrST1a555pLBGPeNo2xXGF7N2QLrRYV+JdHIATgMGCAN22uoCLYFqh2Zg
44Qazo5I5198wAdf3rOT/2LsvVWHgg1pSes1NhQykjVb4vMneYa7FG/ARX+4j2m2
CuCls/Axc0BDu3YPMK/dRhkO3NdUuESR6Bdn9NC+e9Awd3hiYavL4BV8oZx/Ar0E
ZZYn5VJobxyfd38k+kRWQ+uNwYIIIauex9yKXH0ByA1fIhEOXrOJr9vWn80Y9P1C
k6tN7fNKar28Ng8Jzlnc+8gL2dWcM0TuB44JNA2l0vDM9lPqKoqfUBxUe/OB2Gza
yNeQ+rVZj4RQruZO3LS4xzWTL/yCnE15+HpGuoZrrEewiw6N5P5CO3+XnRzmSpvm
USho3TKOTR5bRKQa1wNVf1Ox/Bt9p/JtmMnLvlcoLThHIGP4akjSB/Nimit9kKpY
Pq8h6RMkXSjrJiCHi8qvQHyA0cpjt3Ihn1ej0VUgTZZGkL1YITJS+SXsyh09JR4X
aNMz5Tf0iuAchNfkm3aEIFbQdZyUOmfQDPGgVQY09Xl6wnplceb534w20CjbJ8rf
q1gFa20ZDHsjobDL37daMr5BdMnk1h/OSNqcLtageE3bBGMcfD/uGV/hfzSloTB9
d43bNEvME8XLCcaDzKFy4BodIy3YpnRdBp0kc4br6kNpfd2c4QnUnRa7SI/UHJNk
M/ToQpmCKqfNnNfy1faUzvszE9jbLGmknIGG64pd4WHGHCUagAFyfWf3HXASTYsh
G3OhTDJqbpVMJxENZ7G9ixoZB0RT211bPcyDKsmPoA/TRzFGLJTi0BccWJyHpDmL
HsHClpYoT+I1K23dKYXe72L8J+fhA0CZhpgr1HFBedcrYc44sETv3nDctrmTSC0A
bOTPPZTQ4vS88WA8AzzDzoPHEoOlwFRK8UE1ylREueR10muWsHn/5k8Ub0xnK4mi
Fe//CHstQt+7VkUXQ7YOiGbTPEXZ5q5t/e04zfsCR7FcD75QRLgKVTtJyfi6xdo1
0kIvY14MnZ6Bf73kCNNJVjIxclgW8BGJiPlbwBYpuUOgI0Rri4z5EcYteMClxT1y
d3wOMVWqr7FMpBVJdr63+BtyU915Co+dgjbMQJcF6w1SRzKJ6YhiMiAffa9LmAFz
ufgSA66FA/H2qSXIKJy3gdnaiC0skERpYDXubOGqJCw+oKUPAop0HPwy4+nRUe5l
8aKJwruzSl1a9K4cmCQYa7CIPKLum/UIk4rg3Yuq4U5Y04XQHDqs18v0tKP47Ip3
RpT/rrnacY8KCWPHMiEpk1uTt0n3aVlEAAOan2apCXX4ye3gUT39E03cUurxt7RI
FBn8+rzJbgN3wl6pU/XNbB9W2eR0g/DoQat7HMlC0OSGzYDVFVDNqiJZBO5QJpP6
LdIEl5HzcYiUAHBpoILPQuTunnNuwXT1c1gJGgxPOv3HN+M3300UK0LXDuRGESaf
rGQUDY+XB3BDxJtNaa1x0Zqzvm3vdYXgXbnT5LyK/pVsiMfMfnjKlcq2X137Qj8B
r9q89ex6Ky67H2ARR4tDvLV+7+zMnintEnoz+doLrKdJC7uMTx+QDOjBRAX6nLUf
LxBh13t2bcc++b6A0AuTGk7lTonoJ+1p0osrdk+onQDNLPij2aMCAQlg5fWZWOR8
bkOq82UheWrVg/gG/brQL2WSYTMN1VDkETYlvFkvbvRBwLBpx9syv2I7ejAIMr4Y
ehfl7thQxHw3kLYvOYeLWLb0KYaPPCs1fIOhjBF/BXAMr6v6gTtPIzwGZV5OsqB2
cPwv40SwMI+5pnln7RSJVtDG1MafraA1Z3nqsImeQHXCQvS7K1ckx0BhyWK7wm+r
/BukRXD8trBg5UBQnhbpp05lD6+VDDR15nBWXb+GswdFnZj807T+/mirxzVPOUuM
l/SmBM7xmVSnsdNW5o1gxtlHxW5tNyowuwsAOz54ZauGzLdIGKEPEh+QYTTx0TwY
NG2BqgUS4ydjGFU6ShojQXPPfD7FTkRKdOZggH5ahOX43y9Jy2AfKH7NHw1p/G/1
TNFgbL2D2WTTI1RymH5r+K44eXikvppFUAUN4W6WEKHsXPAsfJDLaMGbFHgg6vck
oWJ4/QFR7+CjPN4obeFTwZ/DbS+RPKlRvJhgdF8YfsPEjCkhAjLesF233dNKplLh
k1FfgVWxwI01N/Vb6sugJz+ztViQeF0TNl4jFHyT2bFDyh7OL/EFq+Kn9aUoap0h
3TQNwcUZQeL/8ZkM45712quHt1hKYEt4meBAu83iLrpWRTI6Sd0BgCnij+CIOeWh
WYShknSoDqBSSyKL6vqht7CqpuLCmF/UDq8pYgDBGd8tmHeKDCvlydOtqAc21t/E
hzCw5WdQZMcOXMcLI8IA9Z18iKROd+13ZUPIjiqaNF5Sbgdn1I602x4AYhJ/kSXz
qW9E4CqI5v34YBQdiL/VnDb+7LheGoAYniGxTJkzkYVKL/FyCG1ugG681o4qnXpb
OEzd8pdNl9pU9uHUV9zbS8VjrFlMWhNJgeW2KNFJZjR5Z7uMdC6hAqTmtkkErioL
7ZXwRhUilCa4fYngx9lLR6b0urk1cXn0sgZ+HQnTHLVh2SDOReNG90cHbayvfrTd
T/v+yAuEuiyztPATddBL3BdqmlAeewztMfff9N4rFKjWAp9cyzPDC1+CgjwgBbfD
XKnjczkyILjciKUhbeT3HEaLhWUUNqPVm636nEPZOPEAfqgDuCi9aNCR6zDhMb4Y
qWwiDCk25u1n7adzjS7D7HhPjTNGslYbfN/zcTN0RacRUFU2QSbd2fbuq1EtCsWL
FbbvPy0ibT4sAaaD2YG2KYpgl1uvU1lWmH3n75G5qd9UfqlYzE+nWKWPHEX/CZQz
r/vDn632E7U0emAIWfwpw/JX1Jbr3/A5tb3VO2Al4xgdXL8DuqRKHlFc1/h0fRZ6
B/vaXAgYfqnj7I97zvgudkOiPaIqbxHO8RoXbzqgoATSSoJCUXhSrEmSFCwEh8yr
I6JUH4OK8Lt0PfXUhWzaE4POTIn5rKpqGZKVxqbRZzhVaaCF5nus95LokmChO4t4
U/W95aY7bhCz9Mlc1VW4cX+rS+r3rz0VR6VQBH2kChsbSIeamDSxJViz+kaDRpkO
jybzHgkRlhZkiqjLRZ0a+dSYrEAXh+KTFYb+KIFwYdPw+YIBIjgM0jTubECpikXF
keo+5BUK7HrV8Qot1sT2lbaZDakgMhxAFyK00BiWRMnJB+MqGyiRiQ12Cyt8Edlv
IjlsCuF1Gog/kwwDlPMHT/cO5+O9rZHtAjaSE6rQf/q+S5QbaL33TymzC8+sLXLL
E+d4qOdkSouEaRkydY2/mxPDS+2rhXNCaKv8TU0Zn8Vt9NUJOLblmH1tXNLdbsFR
B95UhM5dQNKQfRUoYsoCCjB79DCo7axHibBL10yDvkuf9KEKR3jGONi6DBX7104a
qUSMokcp5RUp1QBPnv5GZ3S1OELSGqfpJ3Wfg8OG8VEl15wdYZ2QXZ5Ado4v/VUw
b1ft5M/e0ikhIbj04PZmPyQiEu3euQ5nOr7nmBGX0TmDY3dvDmmPMS/ZH7NExRgp
ftgG5hBdTYPYqpciW741bBdW/SOc8pON0GLaoozhxmJ1JxdOwyYXSnLRyyy1DwMd
RbvUrQFCvqKxJAL+CvZqf2y788GuNOhSg4igZIdiZcLqNquKND3Si45J4TEtB11I
V3JEAebkeJ+V3h0s7JL5PeCnl5lb/rf5LaAg/1Jb3Xt7/r8Xm3n6ELuL6JD2qn0H
JHXsZY75iYrc187nKWS4TTrmug4Yl9yEUjKwljn7hJfJl6MGPJyhhkyLej5qseLl
7CWOtvAPCBebonykyyoluEEPEag+mfQecTJ3l4OGdMOZYpQWjUz9Ft1EG/TGh6Lu
12N9ZS1ss5oqomnn7yvqLpZmlHAKH58ku68RFsEhCi5tJ69m93BVa4NMPJUsau0R
oyKii6ZQu9gv8qFSoD+bbM8og3sKzYofcUGXIuUqxEHpuKxsyVBc8iWPRActOnE1
WzigI4xIeVdBeg94vJL3c8JWZUGyHz5JvhxbstAEsxmxak/2fO0URJ1Zenlrxm9k
Ll3izJ1UqDMXv9LVp4n0rHkY4eFDjYMeNWfjz0p+/ca1JkLFTm7kcjYFMME3Bxxk
88dmlH5eZVA2lkopfZ5UjjZ2YVTTfMVzBZxUt/WKKLuGWlQyTlBDWfIWlhtaQ06a
htv+b2y4V0m1+KVE3/6NkerhZd+Edk++CdBrU3H/0Rwkas+6Gua8lFuoinAH94il
6HjApnowUz4K4kSlCNYBpg0rjdhy5bPRwQBGquwzPChrmy00egUjcpkAHSPs4gGr
n5nFaBtNIYJw+OHFKJPEDlQ5AZA4fsp/BPqYidAcf2hT1Tt5hwgU1nEsdeJ5fQzv
MCdUTk1Mesn5ixuwkjobJcP0MRluZxJWJfZ1GkYLLOfI7q03Ddu1rhPgfpxha/kf
Cb/97pT/lbKeESm32KrCi3wbxwEzSQRSyHkfPaW9OyGiNMDdS3QKK86nDBhe5/IO
ZxGw5jZMegqlEfRTqDevLssfloYMnHWOO90VZI4CRQnHgpHHNJFmHeTzIktb6d8N
IM7ai+ThZdPalmU1Oy56oRcWDJx4qVAXSoFZyeHoH5Gl5bfnTPFVKzl7LwtsrUgR
hOXuOSRmIfUXCU6j82JogeRD7mn/n8c2Nbl/XHbFIWFq7GQXIri4SdJrLFzoPHCQ
2I8lXN6dF15UKy5FdItx+4HVabAX4RRB5qF+VKsc4NZZl4hKYuqWJ3p4YD16UrU0
bRStp8vTcMEvVnxg6/9YlGTAiwh1oZJs2dPvIpvYn7xVw9gSXJQNJOzmwlEqp7rY
QEN46nIy2LG+GRIb4ME1WYAZ9ybK1ECVyXo9E1ddFp5rNdr/wsSHMiv+Lo0p62kf
vQNPAzYWDUGi8heKdl73VrP4QR/ezkkfKl53lG2rIYU/WwmLahlGPpQam9o7Oquv
kQvxbxkI23Fq9aXdVgTpwoWp2t9ilTfCetnK4OG2B5T/fndghqjp1y8L+hpMV769
7uctbNDFGLouiWohn/x6tIjXjDfPjvJCPW8bFWBPvEVkkVMguH+M4zY9lXVbRCTy
rkr1Tro79PNPewYcaB2WDZK3lVXFoDnGM9V9LuC19sMkYwPs9J2vT61RAkTRuQIf
joE7TiJantSk212nbs6sT/q4RLdH6MfmGnJ3dF6oSObYAwELtkYQKcrhpIFTN+XG
imLTyVyHBNyrmiPC1zZyqm/zESETnmTLBoWec8PW1G9Q3lBWZCRi8tcYlahqS7vG
kc/xbzYH0/mmhqrppTf7/xYM55+0/G0lmf8+mo8OyxBYz7dR+U6o/t6H04Laqu43
ftPiv4K4f2lv0CjK1Yklkm1hKWJr/elBDp0Krxtnhanj3+tQnY+xaV0m51ucFZMr
rQXaxttCL/A/IZ4AjCahatbLm9yBQh/iSnV/xj+Fb7I5IN+aSU3siaQ7C/Zslv0Z
pP9HF3wQbNVOwhtidH7guPajkf4Z/Pt5BOkGvgCOHNuMgEkyciIivDwLUdiwt3iM
Uyl0loMCtX5YAUD02lWtm7r13pfu6BNrl5Y9mUiZIO8PsB8ZPOwK6GoAZAo130/t
n06NhFjJ1uJl3/mbwNwAdG8m3WC+2Xsnvx2Ik82K9atHMTjDtGGA5d8jABCSkPBI
VNSVYqFw0KUe3CcX2dmLzWOMZQrO1OQsbRU3T5umNsvqzGM/oPXQ1ioXG4sxvP+m
7Z/AR9lmGMFw1D8x0N+5yjxCk6RyyAwbrvswWOu3uI6Mzh/3SnlBMspyKVmXySbG
jATFXVF42ovXxkseJmKoz/NvkfIrsaGA3oljSbng/vDkVD5QDGnULRFvfNdjlyzt
v/UilwT02uC3up+f5nsLOC+VtoUhaJkisuZelhOFQJr4QzOMzolyQwNVUpLhdcpj
HqsHb7L2e/xZcpHE/DTKWbUAOzTAy7NjuowwjLWmvO9JXnnbUDQAaoGMozTO7gKg
Q3pKnEXmzPjV8e5gCiYa/U9svmENBjc4Q53oIIRtz+ox2n1PbDzE+HiEOibKzP1q
k8kB8lnvupIXh15a7LKpvwU1S+NddLBlmu6sU8dI8AZBrI2XPM8NAf01aPCsV5N8
LBVdoWQ2+GjakQeg++wpZACHOX/4OReXIMndqmHhhj/mY5Am2iIidEg00d1qTbio
jLOPvwSC1cjxyZQVW0T3YB2y1Z5CR9+hDcJkb2gt1JSrYQXRqU38wEmRALyT2E63
mQN6fIsb0KgyzuqwaRpR/KL0iY/qD29yPwNTi1J9N8MuJg8Pq3BiFUlWL9fYgots
iYHfhno7lH4dsAawz/bkkK6y/kJ/TQt5cR2v7Ui/vlHLJQj9VFEpFEMbtRFGnCHX
oD4CXvrLI/eElOHoCYB7gOs+Y6gBbn0FGDVLNKQV3CkOA9T9I8Z4nEK4PUZHQkQt
BeFKx1p6b8250cnFegYvDLz4ykBfKZ74mUmWky+BK4bRm1pG2UfAQr1bs7zT42mG
mLckM9OPxNhkQyjXfvl7m6XZrbvAxxXHbjQgugmq1qgsZ+l1tzimESUHE9BEBA3b
aliwQzdrjZudzyuv+z6InD0AuMBahJ3NJughGC1QrTf8grsndO0mlGZ/k7QYMm0b
VFVoQ0avnGoZVpK2ZK3ifBA0eVV38el4bGjp0XacbggYAmSP7hpqIxscbLn/ls0B
GHGx5S4eu4jkcCHS/Y6wgWnS+MYvgUbAL91KYIek58uZ68U7XZYgRx+UOmd6zBkV
bsJYmwvOkV6Bgtem18ewK331Ft0TGGvNXqhnLApzV51lQtfCobGsC/uDIpp0Y3W9
epFIf3oSeKZU7rYKq6A7HHT4358uFVJRkT5QvDy1P9TnvJPV18FpIDdWAVCb40uE
zebowkFmUhyLb3/Uxc6C2GfEsXdLoGmlMiBt5i5yRZ7yDvE8qEiHXwPjVCoInvxj
ZYex2ftK3PJ51FSptgLwqXvlpxj72I0ee8OawZWxVKR9+DeJHe2xS9d+vdpnjo2G
FntXwM84CmvX0RrFhN2PHk34HB9kyZwnUgAUJDVZOCzoOMoUpgSqlSrkZp3yosjc
i+p3U5a9b0nMq3V+8HW7mUX/fLB0vKeQNZVoXthG/h8KflYYXod6CQD7Pe7h1njw
jFtQxKcq4YkWGAJp0r678sqZt3r+e7fbDeJioq1JpiJUibwJybRtdAgDsBKC7Opa
H8ZghlV+pGvcAkvpfcYR+pDLsEFEH+pCu9z8D82j6ypnkm3g/GhQuMhexJpmahDo
EJu1UtBQ9aZ/SWBYtb+aDb+kGqxSK6bksMn7pJApAnBm8NK+1TXS63MBydr2OQpS
Aaukby1XJurvUQlXRZsXbFaCyT0jJCYvuPFrE0uTOQ/usc3Lpjp6aZfOF9U2WLpR
9ghuCG2pkyZOsJEQ71XCGyhj96CV5n3rYRW7udO/VLqbfuA/HzdYhxLUUh2Oywfw
UII78BWa9kuY9Q1V+PKDsueS4VVz9qZqypUMCwvwpceblwZ9K8Tk0hB8l0ZkUBCJ
Cs9PjugsSDurRzHZNfD1DFBq/627uLPUrpYp37XcpShy/AAVfxHRdkp5nyfTPJzB
R2WsZCKXJukBAkSM0hFJr6kcOYI8KCPfR+vOy2ymJ6keQW5wGUyXCZQV4zx7efRr
T3pxq2i/rJmtRNc8Lve5kFB0AcCGU8/EutgjLAcOrQLJm5LcJpAOw5qMJaZVPkRE
50zqSQs3uv9EzgIJnAhrc7QIUbrJ+MNDqIySWvvzVmHTx3Qup5i7wc1Pa4gM6T3H
scBvmgjWHYG7anP+LKw9181Eqih/zXODzAT7VCaxbF2OUxbJQGfdNXjI+KewksPZ
wE0RiFu6hUNa0v0op99IXRAnK4oFzdqM8h8QkQ/Fm9jCFf/o2Vn53yL3GGDHsadJ
xlZST5hV9YzlRA7BPQXfQLueitJ5AoDJuJKdTuObCJFja3a61/v94ueqL7C9BhEa
auhSMaplwGvu6+kTLi3AX2FRtWXqMhZ7DPVFr6GxfgkkPCHTO//quBXTLejhLdup
rmpRh32aCDUKUWsGMqySA+2ueMirR6bOPtYqYQfSMqz6KClv6klkLsseOhsYHpnq
tr/D0bI0HwbdY/wvSAaigUAu4hC+EJhR/AcXj9odJCsuM+45ZtpliDa576EEBP1Y
nnPUKxWv30+CmRMxu3zyMXFIyNOqzFv+d0rg6ik6JDJ1gZmL6ffBvqvz1QaJBciF
2morYtwffKlOL15/C58T7VY8LU2vtPaHNrGAu/5Os94Rmo9VqVW4okr604Ot/kDE
nL1r9gfcwWU8Py0iA4snjNcRo1ROkRjUgoiou7L2/l51RA2yV6p9r6h1U1kfjX9k
TKzAZ5TXGzvolqFlITKRYDnW+c3Rucxm9xHRDBJ+gOJ/TuOJwiamHHoqDwxNT4+l
Bm7/9t+lyjbn1gosuBb+bnzHcJ238aD9zA2eo92lHGcmW8e04M07eFOokRAu//aH
n1RA453GhBnlJArS4iUu4Y034Pchik7uk3Q+5PTRVtZ3r+hSkwuqpuSJviE8bAH6
QT/jgMAU8PEi+KHEiB9tP4fJEcrOM0ocCBcGBSD8E1ABszzYxP+EmrBw2nyz7mIp
9uXIWnXR3xIjfNjuxxQbMj8ySvnnmKRinxRk9eF1TZpJeGxFe5rLCS7SpaO5BD1x
sQSGXjnpwoxPFTCJ9vLDm+5xZdqKi6VkAqAS/xMwoCsof1ULh5BfbAiR75FBDIGV
2aYCBm/DQN+m66QO07pV3Qu3HKcD3/NJejCoTC2jlDYx+AAh1SnBiO1r+zj7ZYs8
S6bqZM8vqpf5ctL77nBoW5TLaR52cnDvwNqWnkPxpmwbys1ZG1t/HTTbWgtBPgeJ
9eGLrmAgrxH2bWN2UNtZ6xkNxCf/jbELvjUjgFixELUHR5MEyz7/ODLsWB58UL4F
N2rHmqIpT1wt3OOYic49SQ3WSIviAsW8eutXNzT6D/n9cTAP3dHZmgO8MOUU8o5K
fwutLl5cfLb7ckwFHa3wogAfqk4ZRb3bP4H1xoppbC6I/l9sVPav5+aJZ73ZyWcp
XfuwpJiomu3xZiFLN3ZgfndRxFg9scBr1iwQSdlKBSk5zvHvn+5qOdKanlSnbzH9
rD/17T5o0H7RBIcMqrp+mJeSW5p3FVHq1Rv3HD5Jon49WwcbSg6o4aB6Rs8t0bKY
AUFhHNs4EXk0vTSAyken60ohnxoJcd0b+1FXRwzzH7CYGQFoZUzMsdmybHxkK7f8
mHYkHrX9vNj4ZhcMHQd1GlgRDEEBsKG4n8Pht0mnmadhnXC8Ld2Zw/NciYahydrB
+hFa8yAUWMpuREXizvVEpuF69Zt/xmqjxjoLg8fMRgZW9ILgoL6Ejkf666xcs3Br
FAaf8Mcd4ZLCxd/BLT9xX2VwfWWEpdfKeVePX9Nv/N+HZYeTJJaZ6jwiymwrHeII
9P8bX3miq6D7Pcn9uXARHVMWUCUkPkcJEnRu4x/b5tJ1KNbrV1h11spb4py2FLhQ
1LCZcu8MEF92zVxaGFS9QJF5L1vGB8VL3t2gNLmZXsidhBuY1o2J6O7c3yfz/6YO
Q/ENTepmVfVQo2Jau01p0YciNfk7HqKna8gLcRxfVlIW7bb4hCxCL7TFEbVg/mJh
MOlWph5QIFkbHsET4c7xVHw9YCYnL1IJEG6gCRUJNUJuxCS8VKyQ+dnH1Kza3+k3
+q2HMiUhzrOjWyg2ROuKfpPnyD5C5mStDgoDq6jvjNba31auMy5m4LTOfhx8WvZp
0tzwPsvOPW+NYmuBp2QSTmxasRvAPlHQ6qAuyhT/D//n0EA4TEAJbsMzlfD4JwEs
+q6ZIdDxotUukWBVEv4Lia0mte4Ic6e5LK+RUU5+BXVXElMag1XPJ8K+SpLSYZjs
oRWnyYRShuimbXhqY5Zp8zwXcL0BWAD4JZkoA/NvYAI+qEai7CM7rE2ktFy45onk
miTJZ39/+t0pkgv/zbGn75J7WHfdPSHV9bWLz7pLleeggrJuFftDJ773iCbhvmUl
KyPn8PBmpRE0D1ICZKBevkyPTSTd7AAiI1qDnJlUcYTOoiC4FPKh1PuTh6ugY5pj
o5aWYaJpdBoT35Xu7M3KGIVgO8X0/J148GijoiG+Gwvqsk/3FUWowNBuwfmuwUnr
p/tEXuemp3Qp5IBxfOGTWxHnfOmaTLYj3bjg3kgJKBpz29BCm7l5BRq6CPf/X7rG
UpifpbkFP8FKR8yE7P++yqmLBDEQPRmqYoB3C3PQnKL8vhw+FBLNYlDcxaLZLDw6
NOk0Lqqpvg3zQWpul7KLXih6Z+7g4SGVvU5E2YqrEkNZ4XVs3RWktwcPMYmhtwxg
kDZPdNRmXzAfCUkGBYdy8dlQmLE2Ze4Be63zKj4iTbcq3aY+wkdVuXPHEBIePlwe
3flbCbqhCQH2W5tJFhTHw3g0Rh+yDJjFUf+YAnPS0NqjGwAUjH+2oomd0PJF6l3Q
R3y0JLeRJyz4O76glkRWtUbYzDI6kQtDg+yskJLeSCalfPfoaJnZXXRxE/wXIU/W
PtIJ8zGL/E4Gw3NwkNEysBmStkIVw3agqQhMAlf3RBDg0wptR8RECrFSnpPCMXMa
6pWBGJCuXnTOgaInv6nLSUDiokYOotHm5y2si2o/yzEIiHkVORD+kz7j+iQH8Is0
G4kciKLLZa1NbZoC/A+x9x6QJpzT0eVuGaDh9NzVBvNZK/E6cIbjk6jCS0FrQXQ+
rsaKYUX+YUv7ovdQmeSLQeiWzLO2/MqIRT6qK7Z9+5iYrO+GZTF6ANqqZFUZmxWq
ZqAgC6zFUSPV9x2e2ZF9vt+XRNOIMSFnX0yV0qMF6cEJRzaFp/8BfC+H6JOSI/o9
cpC5e8pkCbv2kVi1skn6eZ7R+1ykN9JLRNNzcj8/N2pxPG/5RoSa52ZpFTVxLXig
iNBYM6qaigQ0MA7jUM1D+O4sTxMRitweNI/4/RPHpgt1g2LCD20g8LkZ/go6w1jv
TFS3udQxcfoTkLxhm0uSvywHg18JMonh0HZDrRJRW91AbLzNM+WIc1dLiauqd1Mp
Lbx/ZES19LLaj7iP78DWb6et16EiYKYoZfiBqVYOmVAWuJiNmezuwc6ovHsLPn+l
0JJ0c8z/LWalgHl8bP1jKUQuplnsbbDBXsNelBwoUXv85g0PdcotEVLelC0nkXV5
ixJ2d6LlJ/uZP88iSdUmWeRiiffmSSscWNspKISDgjC74J90KsZUQzBQQX1o7Yag
7lcxRqhO3fswN3og6nP2kWppKi3+vCDEKHSUtNqA5x0WMiHvcjFGCQmStatAds7D
+97KR4VBupsSIL798lCaHHJnT88o1N/hoFqhuI8565awEPmH8xCvpGYcRgSdOM4q
7Fpy8t74FdvoLSmAjzsOjazwESIX4rpwSezeWkl9e+J8qf476D1RcA/ATS8ZJw6K
P1Zsjy05aWdZ6xhPBcXH/Og3eElGi9HAbxluwgxSZ6knbUXaN8mpfyfigJ9yToF4
dcX6PfzMhD5lB1OVS+tzvq5LHZmHsfo3reNKIZkB0I3MJC/CZvZVDTyM4KHq3LZd
NDX66Gc/7xVagxBvWeQA2nwYwIPkBGeq74FLHa7n97OjwxlBw4rYFkcrgBXfjTgD
r2RsSRyIQsLRu8OGi+Cwre0DHbYiPhYzEznvYS0wpY5JUruXTwTwE2frbXZlwrK/
qgFIgpuBFATPXHi3oltPxKROLYXHiN4xdX+2Z0kOosn+RRcuobNXdCaoeJJULlfs
/EBH5VBuS1UkygqNAperNZ223XDuK0XvQdz9cUrzsxc2f3qgk3Tt0nPKNVJ1cw5c
FxHBYztT37EilAzGEHjtaBUz/iY7Z0cngpCV2HAxgGAMzF5h8frSi67GqriqHLed
O1ikINCR/CdWLjtkBpSoZ/8fIf+vDcklYudAND6z5GAoapi0MdtPHu4/DIL8P/BL
WCTPRfgfMSvYSsEZju1QU6ylHxtpZUJiCYVlGubq8aeNzygzK1DplMA3kv977VBJ
J8SDoQywoi0lEVI31ungkm9rU1PBaWcFl16Wo46zHMACA5JGm+VqSmcMr3RXg9m2
ZCMFFwE2q4SifJ5SjZ8+JLCz8JrRSEfw2vCU/giBhE6VWXbITdJzIPD9CVE5+0wq
TTtLaINTgjlAyyj4iu188f/WrxtrGLxJEm4ErJ7aSCMHHmxKhoUlFtKgVdwFcarF
d5HmFV/iX6ch4B5dPNjJd0dKw2D1j3tnumfFN7avg6rFur88+gi7je2p7/rkyesH
dbp9FVuyxPOXnftTbaUb/a2y5hw8sO9SbANvBNTAZ5AazDYvok/9rWZDKeiXTZOr
ndqPxTfHWNYC6KZ4qUAV+gj0KWv9B2YWn0vqS/HHhKuTb8gt4kPWaBhOeytftBoh
If5r42Zj/c1EVoyXG9QLviN9FaGIMWWQpMEbw1NSsbm3gHrAvKKmrhhyWbBv9TxW
7czZlEAQ2i4CdCtHwalIW7NSRYQhXT6/e5gvM5iFJwk36d17C7updy97utW/EO4p
bAHrbel4NUug07i1Or7NBit5wulQ3v9KxR37w7aJtkq19zSQMq6m3+cXBt/2/fYr
QkjT3fuA3WIxdOKa9Lvz6XKM72ya7EU/h7eCntAFx38yS5CP76jqr4x6WDm/Y2Cr
XmAtfLZGsVn0tJUAJP8UtZ27t/YX8cphaFRjN7TCmEeIFY7Hiygfk+YPaPhYocoN
I7BTMuMftFvDUKf8AtNq1cvTub2eI3IkDNGYNPk6Sqyoty1aq0kqFuzWjMsktRO1
XpkMi20bJa4ac8vOX/dygzqOiWfA18CIlR1+Y/hwndy6u/8pNMekPdhJqfgrbhiy
ebx4Se4WVyqq+stE7YvtRVCejuGL1nr9gu1WsjNHR3tQINnSNcG/bQm0lLb0SZF+
fMzXGrMnAHkW4mFhbib5ZejGYTwsXFGH1KVBMUTYeSnlj6gTUmkRGqLKDOnjajef
se964aME2Y0c1qjBI/1Y9JcA5Q2kqQnTcQqWiVpOfEFW1faCqkgNsEcxut8GPHN2
3Ih3R1sFROonpckX1RblUMTEkPu8J8PsTjVfuVqEzyv+OjWKvyfUPoKAqx1c+/ux
eeSsUp+0lVRrcPiN5Y8nOEh89rUz5foO1xPZi9RsEdbALg9J/VrDEvk8nc0mDDxr
av5D+znV0q3FTos6/z1IdsEy9GAp73OG5QM9s7J8T4scgkcJhF4x9H7WVKTbiZ1B
z3Xfqq7FNMI7LPlkdi3BmxPjwgrN1DNfrteL9p5H4pyeWVmTL3Ox14U9BphUe4qD
XTCvpX+GwBuZfnfydcaJrGdsult2Y1KBF7LPcSN6pvMt/rKXxXEg2gGikgFfcjmJ
MUjgoLVHXF+sCztVfMyNYhigY0+Oh6NikbYHvu42mdw5AdpvqjAVjYXv7xZ4KIYS
fBU+lSfG6Qs0PTSghHlCQAZ7VSuh429VKinXys56I5lgh13DEzvXPTHpMhhr0EHV
z/B4GAIFz+sUhKdtcepW2dLtxASccCKeKcmai/0qgWOLOqcbW1p4T0PpjXwLw/mj
H2VYkSi065fZoQxPEyXH2V/ZKwF5bb/+rQk51+8057hW818/RyUFki6svObVJsF5
26cwB5VCErMR2hRv5tEUde9nTzVzEqfmgf3P4fBwhETloNLZrhdgLqr7f2ga/vcH
gn1YC+uPrL4aGfADQGasaRq86KKOO/MfYphdtPxPFJzTAOwjsUr4lEskKdWnQ1x2
7xT2wZusgWDMzDg1pejeRGYFs8WQNHCus+ZezptLAhq5oV63GxPaQ2tR5jP93s+T
Sr9Lbf5ZTquGy+duYCam/aJw4v82g8Ep9bVn0vh/l1xsD0uj4Tc17i+rRqVP+vMH
5AouOH7An7nnuZw4uYfT3pWg5p90IGshjcZd1fEOzCYucH+LXH839Wz89UgOP62i
VrZsBFMCylwvn6i/AkodgAy3ulKy4uGU/gX1iEI8mWcxgl2dhHdAK5kvnhT4Da5M
efIRdmsel5u8MXuesrmuPCU3W5i7oepLFFnFg5QC2fPEfdPBwYPRHb7TOSke/aZI
mLLjz7ooj0GCEtUMCd1teotixSmHj916xVovnToZfkH/Gs551RRXlMi4oCRU/IZ5
7DuQALFJ380NdkO69ak+UwqQTJR9RLsW8LW4VG9F60i1+FL2b1zyEIS6B7z+rDe7
fKE/7GRPQg5SpkfrYO4MJBOad4mtpJTjBpqdkg9Bpw6sdj4VOXIX/JVF9FvOCnnC
zG8ajTxOsx8/En/GTVFbbrEiP5IykeOgnXqCgzPBWvWYrLYigOx2dGNlP/oFtA2o
MCHhbSgoQ20o8DlDDdRKzW6otgSdibL6fnC0lN7YNhsYmeqdVn3NqG5ZJ/MVm+2Q
rwlJ9l8Iu77bqaBfQzQGlE6W1QMmHM9CqS/S4yxjI/WfN4vsJPK4SIFWVHGyriPO
cs0Po4UlA49dxowZUL4JMRV/FP5/avSL3pw+hLlCrha0LFpfaF4NgLmEDwy1V0jT
1Pemacirn8WladkvjxXYs7teWtZcFtDCn+u6E1ugzWj1LoDP9RIS3AtSHq7B3J/r
b2khKUmcxck1bA51h4I/eA2PLNTHLJhQgYGnr5sw3SdxA82BgH74WrXO8kj5Vmex
DZ8Nu6PCDf4/5a+wijEwbwYyN0uibd8A8TuYNnpAGdc78dXvgmaScSRM+4L+UIJh
Y3xYrI0yv5uQYtttWP1n9itAg07nS2xuP4pOMyoEYlbHxaixRz+eBhpNgyzzvFnt
qx5GlMLOMZQdLmnqG9Xz+7lvRfftJfFucZEEfw7G7U9B9kTZofMWRjlzhWjiRjn+
JG/BuN2L4CYY+PZQ80o+3bLbjFJWFtC5frk9mfWUqYGP0GulKGm88NazQVTAZXLs
4+xcyn6SUZf85YFzMJ5PJP7rUNGDRG/MYj6h6olve/ntdtxnH819118CywmXke93
io0LSsNFc1hZ/RQK0mpwuIPd9/FvngEacSXxyrvUDZdmu74PwgxwZeTqQ/RN8H7a
R+gf5E0ltSWvmresbGucf8+0NjB2x2ltwdSO1wquE9CRds+lyudOUeXTfGUSXG7V
pDlVR26q/c7b/bVuC8FYfCkos6HEmMFk1ebM2qmWJfHkfaI2fvv2vUpSBIero81h
5O7D8HSCLRL82NfWQbmjFXxbsv3Vw1RYAFWzEQb+1Z+RQnmJcVPBUcGfd3OsUNom
S1PRxwVGMTKIo9YmLRWK/E74SBbOE33x9yegFrnKf9sO3neGizVEHGnyOgKEmHIx
cwZexSqQTjmUXemQHWN0tlB9cfTjxQscpU3zjMvrPemt8DsT7GnJ4aYBQwCP4nUb
vUMWNNaDAOTo5J3cYRJrAJwMY/gjnQN81wXVnrFq9JHXeBa7lW27KKGN1HRpSa+j
ehWeMYay6czt8AgOQIIsqX3UlkEs7aOIZolqn8NQYPdthsZhYTEfm1QHS1JFd5gt
/IoR7fk1IEA2draBKyJXTw5RXtlJlQ3AZSomJWRZc/rjzURohLmZVamOMX8iSuje
1yVpVwQ/yTvgz6kFKWJs4n4gohCycAEPkIKKivNsLXzowntRLjXjnhCvBzhU4sQJ
OIedhg2Wu2AwFr5JNME2wSbj8BQurrCG5Ujgh6YSxjJ3We+5X/tcAuj/o6Fq00f5
pgyGVkKGS9RkJZ3rZET0hH6ZHGT4nfO0Q2QKEiihsjwa6TAXgQNJrTuTFRHCDCjx
FKRw6OiNJo73Sw5pP+eSWT0gqL3Wl2jTmzjXbZ7O7+1LpqueKMSEgBG9p/C0Bl+B
/t7u0vzqbjqesrZB950vwDV0kToEAfCiKINYYVtaf8TH/a3q9q1TH29FZMIFcZNe
wOBSjycthzEqXN/zMBRrFp0YER+/fzoDQK21uez052e0M8Th6Vqi1mfmBJ/d5bMk
E1UB+MjSS++Vhyz5W+OwzqZUO6boQQk035ekVx7ggJOrcqAMOjt01ccZlHR0g1+u
k231DYuFmA/krm9V18/BEaQU8JZgYkCkBfE+gEVtKrRAWFOIaFTusEMGOmpHlJaL
jg2TlnGNTceb58NxHBUk2bwge59WWmz6oiRCDTZ38gPH2edDmi/T1Ja4rxTO4PqB
HHRbBW0oV/YR58jNg4ph4C/rTJDASAUw5+n07xKM4jUz3ANQX/c17ZNpcqar6FMG
wy/ZpdLj5oyql6huCEIiLz8K8nqH7elEDHT01w5IBI8phZ+rCrf5rcjVYnam67TG
WwaXRk8gbF+D8u7jnBn6MkV1wGdQc/fcvEqmS2jVk7wc+aWY3lDuKDOfKGyRoQbI
t8t43nW0je/ySg65kgdEGdsE9ym6jxQccttFWeoXWEyDQD1hDPX5n/PvJtuw0LQf
GlYxqIKb8jYRBdHwNwyJYmsyJr5+rQw91Su5e2Ekq8gz6zyCqJwFdh6NRmOBA3hv
3M0bmy7m0mOKhVeIyS5aeye418Wd0hy4QP+CIBRjYEkU9yN/Y2HCs0wNe3RSBjM6
J4ye+c2gfsLMtUWJn9vjfv6r9ZaBJJjxWamB+YvQ1JbMG3dXkN9BsC7yTGo2DMjK
p/Mi0HHMfOl8rAXQZKoS19btLo2zuxKD6H5OiLRczjOEPcztASfOYJ1EsC1vtqSi
XyNfgweJWijIrCTK3qWLmBsj9/PsLAgxnoCDuBCEI9Pf3EA/I0dTnkty1MyGO9Oi
0sbfXtrrlsWnqCxhw9/cUDwBr52fcCBVXyPnFdtcSueZEcIbvP4GRwDkmmtUEYN8
W44xbwavGaOMaobpwVKJFQG0akH2Z8p3Qp5hBln1LX2s7Zl97QC9pG/OrVALT2eM
/UL4Jobr1f6ze3GnJCCxPthFYgMZO+KO840ibkHlvaSSqzhhIOkeFA6FOIGzcUEc
wIXXu8PaoqxUAJDaMfjTrXNl27b47sHXRcvOA15VFmTBxkotbc7d/I1EQDn2Xb57
wBsW2IMe3G0i6lcwS47xbPA9MVITKOlBGlLpUtzAdXnvgECPLxSCGQknXJTaKJ4Z
zA7QL/lEAPLVD/5fmewrErrXmcQIBMyTfwX6fYoRL3t+RlKsMDxpJ0QevLvqclMd
yYEwnKGPrlbObUyTGyhLGACBNIc52K2zeWGVn7H9AQHk/GKwKZGcvh4JAeRPTfsY
K/E2KjypqsOCVCdmN7jrIbNP57tuWlz0lZMxx16XwAbNue0dgCNE/itifd/dDu4C
FQfwdzV2o06wjBjFqOhe9WCzVMgepLPomnBMLVZnH5QCpujZJNmeNsZZmhWTYmbK
D+98qPIxkmG0p4m81Mq4OwX+au4ef3+/Kma6If7H26S6ViMTVHMonmOQiEVXIdLV
q27FpjEVH0dXL3jXFS+P6/W5JTGJVwhnHKMTGVmTtpqO6iqyZTBkkpFgtn9HfoWb
Q2/bM0+D99JB0+6M2b2alWC+9fbtI5KT3eQnCAH2RteIivvrIt/LDBAWrqoAZ9iC
g7n/nOSDEoNbGmEfpwZukhy17k9Ot9HnEa8GJ6f2X/GKMZDIBKdZ7dxXysQwhGqK
+DU3ci2Br+QjoVG53wiyrrQ18yixa8t0lTnlvV8PX5pGaAIxPKObkjovvG9XSZzc
jt8GQ5mq+WLnVCWHSmsj9EOIOsxRpIbv59a4HMrg5MgFDNbjw2UCjzdi5IloUAyG
Vci3X3MMbO8/ek0SUK4XLSo3VWWbepQs6eooQ55nSZjF55M7SxQQJcAUmv4NbPus
ALtxMLIUE+/+UN64BWeVJG80fK9U2tGpRtOu6H9q6wdeU5EtDzkd7tZ5IxjOQoCE
Uyg8XfGTrkM55KAj0FfzUme1XB4DDQLOn++ZLbTNiZ0d2PWfp1cnjrBjkPmv8bB1
5rvXL6zDM35gU33FBd36T0Sh/kYhr76+F86L3EwJzd3SZ8ExWeSWvgbCRJ+0N4Wb
3EhFKumss4X9SPvnc5ZuXHChpgUtE8uDlBK7n1bD1acSo0B07M6vjuPR7UGx+O9D
Z4gxcXIcT931TAkG5shkudXiFdQ34fUpxTm4pmrUaDb7A4sKfXSBnnfQlwvxarI+
e4o9gunpI85IKKhZcInl5zD0gxtsKpmlUk1RzEK50/DxaZoEYg1VHCLzTNLs9YBA
tEfLWDI1bbnDR7j+SxGUhkKlIC5KjyBSg8uXFjGK4151Hn4d8nLjIl+DwipC9AsQ
rVO2y/gT37qBiukzGpitOns+usoGHExr8j18c73mdOxKck2MSn1j9txbVWJxWLM4
wW6bIjT1jRUPOBIdSGomeaRMIuUDMEKCLMsqPqB14u4ENfP4DeuxD53Jpw5Iff4m
a8/Iv00Hvoo7VhA8m3ZIfdNjSfNxdUMA+kjdTfRaqWdNpW5NQbpng1EzcXDxXMyu
NoiiX8etMHGXtEGAFN5qrr9QcBj7WJNV/seu/kS00HePEHqJoe7dQABgrP5ekGkG
VgSPOIp0NojCTRUFQ5ghCNsxDV2M2xwaacimL8hSqLB4Ndu0zOMHoO4ojkI2kPIX
rUpihmr3QfTSfxZOw1ctoH60kCBTpKIn3NSkXiJD6zm+uybXB3wGU3oW/mX/dMDa
PkmaKkYsUT1SWloXixPfjiG2eJ+ghsjA88WPyCdEmrzXXuW3hJ5qfPEP+Js+ZQm0
aIEyI3L3PGZm6Na/Hx4JTgeJnqu0Vwi0bSEniV7StoSkYjjbSIJYAdpcOq5HQw2u
g7NhgfagmupMFh4Z3tjIJs6dEOT8TopFjBf4g4x78Sk012vydru122Ymzu6sd4Ws
243suOhawWyV9TgmZKaSv5qFru4e3TS1BuYbNdr+ngwq0lhNq/oNWJUqZYpZcZzm
ZZA6XW6RB3LubLM7CqzBoqKMWIXHsLe1s4Y07t7d/n8sLv8+xiu7yjMslJf7tNKY
ohscpZP26S+FmGKhpGOks/W8vDkOS90WN0jWhpv4CZg6NArkSDaSwGUTGmIL61dk
091V/zVe1hU39saA5heDTbHMOJ8MNfeJyS+96QkxzTTY7KWcKUNl4CUcfR8F6OYE
e27h9PXAvvOak2jTZmqdT8NgRWXPeXWK1Ghez0/t0Sr4jdOywj/8zdQsWY5uYe2M
mc/KRrot8Uz3+1Xyx1fy7ZUBP7wA0Lye/UB/LNpl5eDSuCRf2y4Ss9hidv+hbSc2
nR55gf5vRFE/HwdtcaeC6qB1bIg6QqMmz+HT3EHJsfYMJoKp9j5loh/2UQ2R/FfH
JTX6IbMJF7K2ZRfKOh5MuEkuzmilH3ofPu4vHXA+UIYmoFMI005FaOyvMeK0GQwZ
4cNb1VAl5ar5F5kDlFbzhkxROnMOxk1sJfijLFSoLT6YkRCjeIe8rY9VqHzyJRJs
qYE1C9oCZYXhx9m1hcYrZA==
//pragma protect end_data_block
//pragma protect digest_block
N9wTrvv9LQs+/ijQ1ENHUOmJSaA=
//pragma protect end_digest_block
//pragma protect end_protected
