// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
AhVIB6flfn1U4h+0BQeh6Biwxg+gD1zlH0VGz10IDsj2M/sAD8Iiuvap2y0PD6XXhruREfqxQSu0
NiIVsjdR3LInCMPo+xd2y4DPghzoKUEOSxSB1utKt7mGdMozlwGHguGETfRYzj/RXu+4zkwX6ois
P8RW9GK0ku7cnZWsa1RMfh+bb+e4+EfbDlmPM+vfNFgT9+nM9hk34ORPcfmEHArdBERe6CMHDD1c
Y4ORf8p9hDT6AN1H56iAN6ZCY9eLNSkxi8DzWOeKCt/NM2dFElvSN58Gqb3LdXNzX3lpTXo43yfu
gSZ8h7KhCyFNvreR3aYiJn6ONF2cFscTOe/HrA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 1936)
TkSXf7TzDkW36yFQ3/CgWwgEA2BBJiBKBT4aFxHxjuwB2YjghgGYoXOlLqZP+WgXpNCnoorHgi7T
Uf0pe+0ztVZ/Zi2s9VP+X9NVuiucx9zdwEtvZTmaMwkRLBp7x9rHMPBI+AtImsn81XsEUjWIJD60
O8zifesma0IPLIt7R9/Rui8WYTzPvE7l8yWm66SpxT3qKkdG7a6n3t925VaVV6S+HUbHEcc48eXf
8i5RMtzjjO16PFzHp5GwpVD86VV9jw5ZKyrWUu4/Yo1rTK1bLSIVyI1og2yXnR8fWQpMhwCeI/qx
RnOW8GgU4bpEZsI05MT4McK7IsjTvig11/N7rOzLY/GPnbEA4my4kDGW7PL/6NbDM2f8lMNCugUT
vGWbYNGB1yJnROMRZ6UXWGTy4plIV55zqLIGUGNUug7+U2TEIxgR2ypVMV7lVg9BzDAZdmFA7zGa
ONY64T53DkWlu4s57ExUmYQtlLZ39aeKp4T2HZ4QQDbtJvtp8re1IbJHlJlqSTYyRVBwRJeK9UdZ
EXIrQnvZ1ycLg47C2K52ZFfF7+gtOhfNyhX9BRHdZjzJBO5Wlt69SprH0XQ1wH34b2wtYd3TJ5Zk
sF39vCrVu1JkQHljfUBiQRKoxfubLk/HgtTPEADlbMBi+f1A/hrARhOiV3WqH9/vP3Hw+8SY+Xck
wSGjvjs9W6Bs4HTeDjsa84aDG8mHfYD0as4PNuZymyCBPRRzv0qxwqj1LARdki7lpssbnxFkg2Ei
HYwlzWWLAgPW9uq1t9xQ9db6EoNm2946uqgpdrAwILf3cj3DUgjnrle+IqGCeNpHO5if7gmdAtgT
PlJQWBCX1oZ4opUA8ueF2OOYgi1FsX0znya1LcZkpNAK8U1LMa8UQ+htUrSX8bHQiJLFxuyTZViq
mHenqZxtTtxa2Y8p8kGswj/EHf/grQAlkElRdMEMP21mk1OfnO2+6tQwSKH6hT2XcZrCSS3YfqWF
oQChiUKQFk00sWK6Z6Ki8SlbEYFw/Nh//KjKJD0VWaJ/Ib0lxyWSdjSeO7pfs+Ww/6g5XeU9PiI/
69VV4jEp6ICU2nqATxF1IPudbHlQRNtJMQe39vdnfQyI6nY+Wbq5Zi4mroK27luuv8Bl0e8PgWQh
ZhNPl4OWyfuVUgMbdqGr+CURyMm30/SACv1Jfx/DM5sBnF6a1CryjkKrSn3yEqIgojfDGM1VyGZ6
a+NvgXqCdX78MNbkY8+cKRL2o64setgt9fIfFUDGsRpTNzzHaP9tbud2bAqOHhc7FUrDEeEOAD4e
R1Tii7BcdaSusDnQ6VktZtwGE9YqaGWp3nttVrzTAsa65ELesGJlCujZc5JGJIYr1J8tSQEKvQjG
yY3XA+HQF6UoeEkG2cPkgirueiKGb6t8WdqwPPtR+4t/YiMizHU583zjr/Qfy99ToWF55tlEbEki
lcZf2sNQ8kyE8lctlQrr3w2xk9stoTysHB4mnce1H50NcqkzV3tFjOlgGsUNzZvFv8x5BcBZXjyb
/AO2Z5bAqZTQOF2X2VyoJEgIiBFYM1/ZyKimTiLme4COh9GYtsV3BDy8xXeJgRdyDnyS7Rd5Xh72
28SUi70JppVA9TtG1kluhYV+4S3fF+LhiXV/a0BpyCFoUVWTV9p0GW+rVVDj01/Ldt4H5YbzE89f
FxLBXoEEwMIaYUvewMQKwZYOgpkpY4dr9sOUJVSQku6E9SK9JlAHoo53GgcM8FQZAF4xzPOtjDvA
uzoulCXhUYwAxtXsp8vJpJcrFAQM0C+mNmcx3VSeHERi4OfoI9vUftqcQeKzXbS0p3JF3OhlpHuF
VasOxKKpdNMlgNdo2KNray4V74lW70lmpv6zJ4M7xkoA3S+Dc+3KrvSSp8w7Myv6MkdZV+oBtSKG
TtVzSKVTPF0ami5I7rBra1t/E3/z8hEUG1ZXH/Ude+RLMYyIxaZBPv4P4+ZaOoiaGBlw/w2L6OPn
s2k5Aon4XhNCKynmLTub+Tj89ULvdeU+zdJhcCK5R0kL2VUDiN9GHxyEBjMYAWiPzoHoE2pC1ncj
lRdTswh4T+umRdCxT1ctbP6a5ylpRfVlToqXwmX6T0nGSewlqKjF/WSuW0njwIrhcJ9jzCpVphaa
65fN9su4jxpUIpw2A+8oNgmMlCktTRxFeY166t2VHnxG7g262WWexG3yTlMEV9S0gsvpwZiQ0TtP
MCH/RiK+Kvhq+lgImR0ge2bfUSySFIWea847c1HPncrRdfUI7endm2UUWQQcEsFveK1pdbdjeOVa
e3qsRTsVkI+WIwn491+Io1bLaEe/g52DGYeQ7DBbZPMG+meTcSY2g5kHlqUetEkT4RFqic1WDpII
JziYSe18PIzz4pdxq7/DzF5S3YrCX53iQUduwW7sYVGjOZBjGMwDNR98hCP7+azQm6TMKQEAUxyX
2J5frwoJbQK7AslhC2NhXBqXpPNiDT3uptCkv3fu1AuLLIj7mP4ZDVNKV2CyKskXtLQX7hFuz5o4
ZAqKhh4GvRvt/lpX6CjcOIUV1ILcnPE3cJfGqNdktl7j3qWdJ2zg2hs5z701YlR1E8Fz4d6Z5w==
`pragma protect end_protected
