-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
YZQXSdbB+U05HtOXXU6NDGgR4iS72cUPXPDz/fvNgWihNsBD7lT9pjrV15OyWzxn
K8WQ8nJVAWlBo+rqZxk1mTsXDeymyIoRExU6ifjyabsnceye9ZAMirokFA/g9DsR
kyKiEZ4BZRRXA0CNQD9I8JQBLgkoz96GJ+Gj1SLa8EA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 7104)
`protect data_block
2c7HL3t9b3faZGh/SLu8YE+xnvwfEZ4ypnDSuFZ7yBfrA24QNgdAfaZMJ4PCZJ5g
YRlVEeMpOAZXJx/+GAHPui6KLMrkCm6eTnV09Y5/FuKRp+fYg6Zuu5coc5QRkGfH
UUS7Sji8eVQPiwExyWT7PBlgroo/CR1vxfik84tZx7vhZD9+BspOur7qslS7RvrM
KK7DUxze1yFa6uGw6wqvXC7YuaZWdFixlZ5bwIGbk6xoUFjaU7Tu6sYBNnOo5szc
GOD37VKbZPuE3vTtlm1CsNP538sSbo/IN62PsijO8tfj6FUeCzvbNjBjLY+vmkf/
m9ssVRNj1XioMvbKtyQZbDpJp9Bk5OFU39zu5Y3jzcyOO/AXdL6n8wGBh9rfv2WP
0MjZO5EfmCmtT9I/9aqEspRYHYZPGF37WZpzAHb3Y7nESV5icKBR65SqNR0/F73H
awJReDxt95zcvZGZYf8Du/1pU+o2f1A0c9aQ5S3ggyHDhblLUNixO4Jl5i4tGVSa
Bi6OxTISE3kVod33lgV65M9RpF/ukpTj11B2cBuCm7jWjz6Id2Au6uDWDpf49f6n
GgzDL0ZYx2TVfyOd7esd4J8aVtlM6+/lRMMntM4xSghMHmt4Bq+5xIuLSM4pdBDg
2khoMOkb31ohEcB8mZbJAXsDiaL+ixRaWl3QJDkybuGVuuU/HSu8FYa0vx/Nc2Ct
IHmxkV1alBoZFrKG0tnu2luIJkKb2669zzYMqM/QmsAEe9+W52+oFRGl47c90AcW
JpWwcGVJd5YaOON42x54qaYdLmwD+czB+EMEbW6BvjuRCDtFvssdUCzlErxXXByG
hEJ7MTfEuHitn9yxM/Ntd4QCNVAqUpgbDohPxjQSD8qE6V1NJAEj5Gci1P4swvOi
gIzDV4g0bgzJZGEBiCzKL2R88Kf9sEf/iBKMFsuotSFAd/Wj/t33DiCsG76IVRwn
2VP2oOQfXDPwPtnZNmuAmyWCxdAy7rvzOBiZ4fhK/SiEOOgFASFkEBTud8btWWC3
SQpoG/ujkKCLFV33VpFqjiyKYgS3RL2HosVKHBsp4SYsXEuyNMgpvvzf+UPcS1cc
i/PwRwJpYjsWeL1csKB3y2kDUqOIBALcyeKsuOHddh+tfAA4e3RV1+wzZT8wkliu
Ap8srNg/fveonDxRDGSsf8MfkkGkxuPCMagxv3z3nIKZgRAkWgtwXw4cb5BphTD2
DxAvDtAQ0FWkxvirG91IL9FNU96pWQs8zkmY/ivyMApIfEOJOLUPBytkhXlj18OU
IDeGAqp2ptsQC96WYLHTQWC4I0gzyCTs93spLgizQkRspIKY7VEPJdGqLa+1qDQG
2qLwljeOpF4BaRa/UvcOKgAK5JO5Bi9Cj5p6MgZgfUqzWiqKzNFfbRbOtJYWekoI
u0MvynE+tn3iQ394EetZgzQsmxLlOxFaoXV85VYbF9LzfXx0xzS+0olQ4UuLWF/Z
vGC2dN6syiIFHeagBz7jO09SBtER1T6Xg7KDRkRcTMX9txSMXOA0znuuZ96fyoz/
JxuUZuEcw8F90Dr1MWcUJow+mkgG2A/zRY/wDZUhzB62EEjnr02f8WlqLJ21/SZR
8TQo5AJEUhmRRCBjnIPWaBoe8sgjXwzED9mo+bZSVcEVlmHbYwa81OzsRB33qylE
4csOe0INRzZawMO51Ms+RCtxa3lNSNiRMRI+8XR9kofAid1APjp0A5NDPV9fXVx7
IbJdrXsFWvXJsR12ck42MygBI8G9diKKidnUFARzNU/y1GNjTMUBMB5QA6dI4O2B
01hd4ouav00ZMiNEG2uki2k3gqirE2tBw4PxhSBW3wMvpkN7CjgR2hO9BqQxDt9N
WThoMNK1FYCgEFVHaGU3N+WF4lPGlX4zGIjc6xHTwTkMgHZ4MVVm+xiZCUP+k1fG
BuIqqUxSWaz8xFhGn4pzB4luuNprvK+zx8kmZEwbVmcFHaAPnLwP0OoxmLghtc4V
+/F0yTMebulf9Il+IrQEMzEm2jIdAVpm3ED97M66MOXrUCotYXWdVb17Es7rd9K1
tq4uDUeHvBdHU9DSbwyU7jQ1KPnfKsc8PTiD/+HH3D/CjnTCezmZG51WpZ4c8k54
6vexwFfQIcvrKm6+NdoDrJllIn/ZpGjEISVXA93Im4sumygrXNI60i/UBO3mObtY
rIsGNj87P2mLVot1VC3RoeNEgu2ljLkONycLiw7jfMkptzZHZuONs61OZYu/e5bp
RNBhxK4qPtSgAhd52ag4XUOwv8dxMcpFEb7u9lLFdhccWvBZXqntq0KkL1OoFytw
CF+SQNl6pzCjKg+HegrtjRKAjm/MJP8zUfSacbPGW7g8jNehYVzJt9GrlvZLxUJT
GCvv3a0TpwxH0m2l/rHQPXVymLUBZpCu9IPIdjIQ1dNNY9HFasDjkmYoeGYyCFMu
oUktW1y9WjTnGf9fwHI1+/8VK5pDZr2PIeKKjHm/iZktz2NcQKd6N+qlbT3s0aPJ
i96skg78DvxGGIy8Qj1/+KlNIA8JH4EIJish8loZFk/Irhui/Zdo2OtoMQjTG+L6
qCNo3hDe9WcvxeHQTkiXfhdJLzjax+UPDjwcvBHD7xjHrWIolaIrRT4U3PhUGGFF
Nie3KebomAnt+tj+sbtU03THU2IWrt1F63fTUiFR4iLVNo4atT2m+1N1/6m8li/2
BC9EaGeAeH4hE8tTfrAO5Ll+TzI2+Nzk3oyDv0mZ473FO2bwVc+4HHL80vCvaE02
cMrl0Fn+jVA495JRt3Ec88MGp84k1se63QOeFGlB+CS/tplFGHG2HG+auy9GHomD
o1FMnpQQ2y8d5vjA6pWDxZb8UX6l9Jni8GpHlnqqNiFT2TuoFlDisg5yRdVeTknm
kXWwS65GdqedoKdclaPEuB6AFzAiMebDveNwsq8bLJ8HdJ34mrA7Qxett8nG70/R
iWgyCozkomNNSIajCRkXfMwDke8tFLpKA86tL5rEl+ISs5yLU+pJHanOujYEvoKs
/E0VuuBQAUV849ZEs9ji8pkY40jt8StfAnFVxRTjhyy7EwTQlr3mY0qr6VyJjAsp
wi7QGVzHlRkSjIbrqaSnIlewQS0n4FAkKXy2vFqmrCT+5e9WwW8mZiZ9bnQi/EuU
YQqBFH3nGtBaeyzsKDhIAqnt6CxW+4PO/EzXm72gr8LhFAPJDl0hMNJRurGuEt+F
9ZfchKSnlZK0A1Bh6rZWQuRTssT4VQShuzoDNHb9lkEXbgWYpc9zfC+WptfLMIYN
Zh+fBvuHxlg37JIRzEl5BTAevm8wZkNKYk+a7jpendyG3ETAD1VdXW/bsLTsKDkv
Wg/89uJr71/2C2DKFXXEtNolwgWfys9cBPop617TLC4iU1LtSsnrLYUPk34aKdiQ
5Emfe2uso4r2TI5T767hWQ9Q6QVl5GM6dKyy8M3luZmifNRonw0YG5hVCFmfFiIY
ktvWSQKlhyCiNrNfwPBBRMLJYRZSv0GymqguTbZjVR1VdmqDXbn7oPEK8pt/Zjdt
ozH/BXqXryWsRUbsswFEqGRsc+cjn8QW1igLa7+N7r7qzGhJarEn216VMpwBXRQZ
vke+13D9V7xoz0ouCrjpOX+ftbUQXFUaf9/OotUYIeEyi9ljJ6jmXzEUqBXXEbSn
HnkvCaguAwqj1hXbD6AEJ4D6TPQT4LbQRtQK4RuzwGA3ELorufD+w4lTnSiDah1c
JBG+tXTDsduBI9cPzPSDwUY4iLrLtRgUzdRmygcYfaQweiqGgxaXwgRmqwlgBkkN
7GpvjfmNEf1aj1T58TY/Lgd57YHUvdOyhA1mUcXRQE7Zt7g0GSd3fSxbJO+uxm60
OQUwL9MnkgVW41VOoz3jodrL7hQMnHrCa6cpyxi121JpX1Uns/ird/Vp3rqraI85
iaGEwJLZZDylDMkTdDYrymdgi6CkCyQRMOy1ceoAYVCueLGGdkYqoszneE8OUCZJ
3+//yMA8NlN8uIY4oDEzEr0LjFyyyVohC1mTpeVTZYz9BMW+lb5M+3ntCjKtUxiS
QyHeNpPoWkyPmXM/4OwQPGSbLe01w4KrPFafvVZc6LTqYEQ8Fnnj33jWi2hdvQvs
EztI6L1rNGqlJ5tePvEobM6t9btx+3jqQtAE3/xyrI/SKVcZPT6qVWVMp+Ie4CNI
gpG9cL4VGLnFHnES9WvjLClvRlu9bZfZKZGf5TYZuMJYg9fVUURIM7zrpmaeaBex
4TLPFSm75o3P9Q/wfMmD9wnDW/DjOhIkO1kbyzTdou9dCrnkuQjkc2Yv9Buki5Wc
vjzG8DJYYjToCjrDEUsWpq+tseK5eJWLmdVGgh0b69rtTc96mfoXeEH31T1kI/HO
0KlrH0NmRu4NFeUTcXqk2XFiBAjk5n7MGxU+yxIoyUVM2Zfl8yBw5PhyoWLAwcTV
jqLEanJsrdcCb5+CHY5w7XinE2Dpa0kf0nQ460Argr5zija3LJiD6z17XXqnWyGy
+qBYMDp3u7fh9pnEwI34Ca93qIW/4HHJRL7T0LFvDmehlD5ckFV9B54K7pFjRoUY
vYDxjlP1vJI8LY3B3fO/6/Hy+AIx27bA8QndoW4WZ/5mXPiXVxUbpKdP+GIGK0Wd
mschrc0q7u7DGXYj50tkpFWeCxlBkk7TOvbsFql/TcTBLiGXq9m8yWXfKCP0wLbQ
x7w0MRBCx/PxkLSgY1vMhheanzHX6tcwb8Wo2ABNmhmqvtS9iXraTc/sbgT3DNBq
w+5mCiHyBYcghf0aLxOVGXgAlo8gmNPxioLOuZ1HZ0wDDCwuc5n8pitm+zMFOdgZ
aJh55CGirapj+jqdqwG1WaZQpprYrvAMwtGIvsqqnaRNIDwrtDZ38FsdK/84otMh
7QM/vw8g+kNqq7MUjid9tcBtW9Lqo/BVaRvD2ejPA5eog1/xhzW1AqoLoQIlZVlv
IQMX93KkELJtApA4VDte1bEULBcApQgQ74qMfFs44oi5iVwV+oHV3hwJz1o6H/nK
djSJ0PzcI7X1QExRdbBDgWukl3TJu7bDLpEY6xsl6bTFX3p8xCda06V/JyRCYhqU
Psx/RoRxIyIKFJfZxkqc6+IUBw4c0p8f+T17SkQB96ekdsAmt6GQuAhWf/6Ho/w4
iom4uX9z6XFSCW61uaNNnQ3n6FcqvTTphykvORLDxHqo3jU6vXwtwV/o67MdnGHi
huuHh2AzOXvPd1af/FmdvH54TO/JuVOlriVeEz1GzcjlDLnaRymVJhHztSZ+9EOR
4QGHq+JtJXxO57qIt13CYgPZGGnmetRyFan2mDrJe9UrZcYzfNDyBFGNJef0TT8v
qss1wQSMpVL3nfFYZRLNxqgFoaOuExYrEV5x3hRTOcGfkcoZJzGPOpXcrwGSUcKV
tALZZWxSq19zDSBvGgJH56Euv+sF5jLeAT84yxflmkuCn4OIECQVok+NMV4+Miyt
qqtvyKffha3GerodWCsBrdHuX7GAbzcAVuMu1XZUzWQZnHETo64llXPudqLgAO/6
8jd5zxulPAUvqSuhzWlgk+hav3lTymq4A6dp3h063mDNS8EUtVNEx3WY9uTxAcXl
0Ekeor0UfZY/OAAXBXXi2EYYyMHxjYyQbZmfXzmpFGYAxAAr7eLSM/bTK42HrGUu
BFAVRWxGME2QsYt6BBLpeKimM1SSXepaIyJhwJzXgKO8l8UWD83UvinvLufRbjOs
9/JxyXGoan3AcZZTlQGumCPfuBbWovr8lWGvbRUuivB6hvmeG2EVCc+oFR9ztmJ9
+yGjvh9V9cnN4VjzyY43HsgBT9BOfYVPs0UaMpb0AgmpabSevwf6ANaLlvK29OVv
CLF5HW6blZjTZhSV0zfTjhBCP4rKArPp840ysNefefCGyyqxgTOT4cjuhxNAb0lI
XD6nupWwYlR7N7s6wg0tb6Mk4xCt5boefFxWhgL+OBnt6NYpFtPpZwvrHFKbFcAf
p+skszX6jQtUmD5/fyLF5FRRIaZdc5eBy/wiJMZOc8l1Mto6BvBM1vlrVONcMbPu
20F47xROrWYVLyB72R93maFMDcmg7qj53AiUi7zgnhU/BKgE9mKQ+bGzyVGBpMN4
noMoGgsy3jg83Rs61Uk+P/av9+5oEw+4XOKjYIB7PgVd7/qo2WG88VoOlpMrXwwV
6BPJWP9f7DEpnb7tambd0eqiBE2BbGMUBfUR5zBkEVdU7Qrh8k0fryTjY+F9m7l4
/vDebTllekYvBzlm++1QP3ptsKIVROSebEWuFZ/9q8NfUyBL41s8lBnXWgnIgbyw
EijS6OPcQFg3NpAP8UjsuWaS4cnotapRL0tBtxywTKxBL/txb5yNHuZPX/zVjz5c
hsCf7U4+b9RZHbf81jQWuYohMPmkMPLD3Hyc/DgaorIcWn8faZ/5jgpiS57FffGc
k6o4u89gC9TnVFmkgtOe6J1ncNMsXiEuzRb/Ue5Xi6JomUFFfnGHlRM9wpddYkTS
Wt0nX8+6EKzls8Fd7zMEh5zGedVl2TYZvqZO95MPTaQo1jTbU6Om045eCI74eK8l
B7YzA/8NjNho5PKEQuJIiVfnmAktP+PQdZy8UPARdbbxaiXWmxM6U5TF73AaNZmx
UmmCGjNlQlSo7MryBaESharKS3ZRaj47j0TRgSw6Nov19INe1nef0JGvenEbVbhA
dBeIN//PxK3KFO+vVw6BUhUwzJj6RrsIHRYaSrKf7dFEQdLyC4ms8vln80IfERrR
s0IoatA6dY0+ydgh6OQGg9+7tgo6lY40UJjUHD0BlFgOPDbFsTjtiah0rdvblyiO
m89O8Cen4Rd5cBWTTRa6JbUa8pJ3IHUnP4JmTCrrl0H8MHp3oviguZLjpimasiUp
wFJ/lw7cEZCEe3bzE7XdUO5BUvROnIjA2mqRrDDGvEvfaDBIfnayVtoHO4BsQRED
GuCxkcMRLJFoGeNNXqLlm00pqxEL6PZ6fcaN8VEfPRVNCxNkX53D3WGCUjFaLkHW
rnp1CI1NqSzQ2agDNvFGvIGLXCgoyI+4txBkoQT83iMea3xffqyiDgjuHUQce12f
skgIdHuDQdbPIAAPnzbxh6UPPOghiJg8JwmSOSoHpfbK8pQ6S6ItjYAWVqsXdW0J
pr0px/zwfp8VG/nw5iXy0rFoL91UbkZQUbFvZt3HeJEkKv48o8rTRK3xoMzZuxhE
myL8Q/d4NLTRUyXUYjn3pl7xvxFndQbnVNN+KBwf/7RNtdp1Zs8g/u8zBEy+v7PB
Tak2v6Z88LBHsO0g+FiHO3IOfKtHFTxkfE+5f55INe2WpwqIDnS7sdKhmqQxBT+h
xgJJgiX04zYfL4pG6tyUsymWExn47vUhxm6q4UPfXYFDa0Ro1aQyjboeqN2HmDi9
wIHBZ7G5/v0Nw6koy5agi1AcZQ+fNvSXly775s3yHoFh2MBKN4NKobY1teEJ0qML
ZOw7lPcE0cJIJ+ME0rK2YBp5UwHeLoLFyakxS8LJ70slvMaHNBJ49smo++uthFQH
ydNLvor/n2pX2D4yx0L+0LakRkgKnALT+UmnAnFNdxL4MDconMSTGgXxHD0K7eco
gjQZEpT7CV9FeeOFI1O/LIRigsdsSZiwJGChZg6pKyhKQde7ACN6qayoavD4dn5p
Q3HARpagblGe63a/LcmFxUpYN1VZw+W+Jv96s6hFKCoNTqRemTsEmXzn0vp2AFmv
7OQh283Lpol3rDzlX4qglAu4OrM25yqABeNLH3bByf3i4wvSFlp1XnrWHGkZFylB
GhR5YbRJ/YHM1isuRuGiGMF4/6xv9eLLmWhvIOI9DXhtJm1QQLDyrXPfwOE69xpS
gvt8iU8AVYJaoA/295jEZFpQC0fgJgNVd6I1lYQ9PPWD03ux+SK5Gcbdtk5KVWKv
BhlSeUEEf47wd2fpYDnK0Qi789M8QYQ7svwgNTTSq6o58EwDrkaHsH1ydmp/jcuA
QP9560W2LWHHuSiIbGaH9b1nffGQ7VqooWe+VPJILJmgpaVl2+nkGd+9s10AaUcp
8VtCW1YK1b7zGMEC13KOLB8aUiumCGEarGy7shiPGB/mclm1HGZQRXhNXrAfINhy
4Z6tdgo+D9JfHCC8gIwGlqhmZcJi1JYSMaoN+4rSOAv8XEnIKR9qnJme+ur0GV3D
sUiDF8VQC6QHh9ylS/IxpmZPYQ0wm5c884rxBe4Y0SSi8qgwKu8myzVbk9kLmMW9
4JiMGj2GalAZZzArOhhu+shK9fj6SOGGOkTaNXZyfSJpS3tV5S1Y+PWQisGIi+uS
9d1aaDVJbOXbQrH2OR3fWdQzqyJX/891KgVhmbZbigG08459mqkqEgLfek6+n1Mv
Z4FgYWXa48bcdfvCi5/5ktGH9DLEuWo6INKKm4dcydZZWCdkXrLzUFku/9zOe0Zd
KJHD1x0RKLE/aWG1gN85KT+GOU77aFStdrlVZSQQDyyYP+lw/mHlR5Vt4c+QMdFR
imVtrQQi7k/mTSvKDgL4HuOTAC9ZJfS3nrN7QekrnI4YLQohV0uSxPup+HWxL02g
KSiPj2mZJtbvDZd6H2CCg13YfjbSqYSXwdo1o6/WCB+7H80XKo1/Hil9D2yjqYv4
uzQPUcNwyVl6zeYS6T0aU4BJD5aJb4DlZYbGyGWxZeuROuAG1TB6HhemypBAKyD8
ck6nmaRO70oyv0NfVmaC7p26IQTG5qnbQmUJKqkOo0rqtwgxV2HRIz4pqTr41Q/x
xqUYr89Uw8PyHY7L/q+AKV24Y/klGKdagoWapQLcdmMxx0FYIUqLHzM3Kef/PVDM
DvXQpbV+EDZ4OPfoT8GS697t9uYDMQr8AquTrxzmG2gIM6RLi/v4BNo4qkWK1om0
iKfT6bvj+tfjDMfCKb9Sx6YU5LCfkbUBWQ5n7TckL/fEH6hsINLnroTB9PllEz8G
98AQaPjPpYhoLP3iOb+UZ2qNFP6M6c4AJvVFEMCuBQZbL+VHn5M7ofA9PP+GPAK2
x0lR+BHjDrtSGS0KFwNpJmuRTo/72urP3suZtgfxJtpJXxCp2tm54i8TeL2bBF/F
eJCyB0qvkfvrpp13HrnORpbIqDyUqySZ2QY1oMyuWGbQ3PWKUKgueSvi9Q3RWYR7
KWoOXX/9WP5x8Ll/2HA6M0YrjAm5vkHOf7Yc3Wt5ZVjGPc+66iEJmE+/kPKEtKa7
UOdP9h/GlaD9fHOGcLhbfF9VxYaQ0/GaGcatXcCD8k3MKhCWixkKhVlnwrs6FkRl
/GBpXRsi2yj2GNdLea2WTBd0WNtzZT89sPW3qvx1cQbARXAatbL7jODEc7v8CuPU
ROPNrQcykPl+6RZRYUlwUoYFaZUk9tTMZXXx1hjUdoDkdbBnJHvFty5vYvn7StNU
n568em8rjjNVNOvIdliK5m/BBfzYmyl1DCFW5+wdwv+P0kGTTM2rFhl+PjSIHXaO
ty0RNfi1sh6nH69KomipwmWaRKmVv+m2RVHjwjq7CbdIxLnZcxD+9i6bpJzKYEBU
`protect end_protected
