-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
mW//F5zbRjZty9Ry8+6KX5c/5wyWvSrf0cG+RS5+1Bab2QLT4+WAtor0X6mPOB+u
2b8ylvosYKiNr6Wmhd2UwjhgomdTofxzyw125lGQqvXCfYTne/cii63k27tWOydB
XrMqoixpCk6QC62lbfQpBjMPl66Ek4jXhV1rbWtwfyNQfw70roIwEw==
--pragma protect end_key_block
--pragma protect digest_block
AuN6PR4+RsGoWZnp15NPfzE7z6I=
--pragma protect end_digest_block
--pragma protect data_block
x50AQzsT3/ygY1oFwM82Z8K960budkYdG/2j7N061VsKqZ8Xfsx5BKR6zYidhB4J
jPhfvth5HYCryyejTAQ2OCElKaPH22qZEP4nTbATf89vqCZ8EEmIyAEhW/HPhOvv
ic+qqgrxu7UF6VqhYo5Vv5gp8rV7NB+UvIwd1q4nYyW0WRHv4Brrlm9VGxrDGak1
x+rVrR2q+2Utvr7ghI3/YnLD5clRqPUT4xf8maLOdm9IFdPzN23bxBfe0T+tSyQL
+xHkP8YX3YedDBmpoYXWo8xYom89fuknelLV+BINRRa5hutDQfrmvPJ47DCk0SqX
wQu0XTYQTawL63oUZzkWi2FkMhgNF0jBveuRdgoWAGr3kqiYTlN3nOVJOfplRV21
FwbNptpfOb+IraDwTKLgA/Ie8IAx2PV+plrsHKXUkhpS6k/K9MIR/+XbrPsvQq7p
HwMRUFpSfDPVYpj/nXH+AhWoyl8k8BZqqOELY0zbhkSC7MT4qE36Ap3Tktvy3PBl
MOyJtn1Jd/mcVulAVACGOTD7hFwRxb+TU6e/EpQhfNpt7fHiV7jVFANlajdAVTRl
LgaRg9gUJMWuwJV15MEhGZXHHK9RcNswmJRJysYRH5zW5EZK7LcewmJBKkMaV7tn
cI0LGAXN3K6HxYo2bOo27BTeV/drDgokCVVQ5J8YApDsxXjfEoG2cp7D8LJ5eHjG
Q4anq6Jl/sD0Mq8DfY3KKvtwIPAG4sKYtwGfdyCHDttFnIYpiquubKtjENANQgT5
eZ9HLNgTcu+FSeGNFlHAtFQLgrfnkM07DUqpftsIp0kTQphAcodAThNamYdSZVCo
sZrSQqxOe5pmaDw41p3eEUh/RE+UzB6XfVMAlyWHqaUk9CA+kmX7SiNYv3fusyyQ
Q4uYf6NtbRLv0/bxPKIvwrHY7Wslxv7aGy6SJBwnrrOtBPzRJQB2iE/c6EsQOryE
+/HiJ53ctg/qT3aoPbeplAzLjdpev4B1JhHaFk/DhInbFdjHWCTTuTxQNh+5qBe7
bcXR7Cv/Kp/K0ZWChAr/u2m0cgJpza0jL2zVdHnQJyB307fK/MjglQtdYYRyxyZh
ZyTSgQ7AWrE0Dzz3KVqEOwf5cJCUFt7NIsxSd7g1KtbuUyf1OJHA36SAWRT6mrBg
yryYrsEjkc8cQ7Lyy4DVhlaHjsNrt9AGNHTYOSs/FqZEyxSWR5pksXA7H/wSX84N
yddu9Ub9tQDWKvQe85q50Qp1Bapb1ncs2sMlz2u0Gz7nGOuGtrc4ae0pJENxaU4/
VOdTK1wyZW/sb6tM6GEE5aVIQP0HPFV+8qMUvbOP/ZFIOEh9RFp9MzrJl00v0tnj
v3zovaEr8yhYQ2jk2S7oV7VeLP+lkxmafUu/UO2XnucSNB5GUFwKhO1zsI3uKsrd
ffnEaHzt8W0tdKRf4eI2vTOrQOIM+zVqCGlg5jDtseCxIecIvTjwrrc4oTwsR8dX
UviLhNWfnxsNrCHtb6zfEIXdr+SrkvG7TCmUER/AuMUFxa1Bdnugp7HYC8jwlYwm
o5gSothykipFBpZbjbxkrS5yhX61lxWIxAFOtl05o0qXYhabdzkzzwYCVJJmlfPj
44JicphoYwkiXcEGVtBo6xKEqGp7AxBj/qL+/TySumcKdXLuLvGIrJYwzs9+Jbkk
Y2XaBFsdxL7bBu04imj2v5jUfQaQhP0mvGhMWnKmiqeKY+627n9uisbWF2/zv/9X
LzmTPDILSm/bSdTQh2JLDDwA3mXyDuSF9115ZNqHNTK7t607OArmc/XJTdR+y4lJ
3DuWsGQIPmCMuIxsHHBL0Mo0BoVsx8W9z5VWgN+5B6mU+vZv6AeBdpk0FA0BEYRA
vQO1euCOBzacmJPp1EgJfGH3zQSvCWa1Z2XjDTX4fUQx4EzKvPCLs2mNQwPhS2wv
OtEnmX/mXVZsjuFz569O/Ysa0KfkvZce3Ln7e9IWHrM35T/MZ3BBKtTPlGYB5qzp
z09zpE841/9uUlWlFfTNp3SPTxZjkKYg+BGTUneJ2EQPoDW4AV8jPcFh7ZDFMpsD
lGWC42Nd2u+O1SGA+QQ2Ipn2AlEb+eeT57BYv24jKGb7Xzzys3ydEE15ZhiCWaBv
1t37wE0fAPClizD7sFPauTTaoBqF4iJPmHl7RI4ycy1DtzEanqHuUpKEQv0bJMee
gSZc0YrBfNi77jPCZ/AqoSIMF8nBfmYwzc5/Uil0OpMACsKAGX63+MN0vGJ5JLHJ
iBiPWi8VlPHDLZwfalsU2jjVlk57IBP33ccOpOswckvlaVSFYxiLcwqpGfU3pZii
TG2uj3A4o0Px7N0fGjQYQPaEIgFmGbUsnhiRYAdGuhFig0/7H4T0WO042Nxh2egR
QTDXPx4KyLpnbg7xMVIoOTs5JSaYI7WekWHAqzeJt2sZ5tnwoDzKPhEJgGJ8kkmv
fzuNQVHu2IdyBqEyzZQQ0f8scl/ibj9utmxZA8j89b1iArGudSOZTmHVDaNzBjjk
ejF7/t3GWlTdYUOht6JEnrsxGRKEy7kawT/WfOpRNUgcr8pbitujE7EOas+166IE
N6Toio6zKLpLSDBB4R7tXm/jKvjiXmJMrDUOnou3UXypbMMgp+LpS5Ogwv7SboYy
LhxvegiC0H++AhuS2Ev5hM02+X8JPWQZqEkzdICGJ8I8dHJ5Hb1LCB4Qn85/+U9K
6sqwzWySTqSv4S+JNRRwr8sW2nBvfP2jsWuuT2Ykd3iLZCRhGSYby4WQiK6dRO9E
/4y9+z148reG7lwCw5yi5bTPLFfLciANMLW0oQx+cr0f7p6i06OQSUFVc2p9ffRo
TipqsjSjyUqEkKmViaZB0GR1rnx1jWtJeH2zVu7zePpbROBYUKyhJ31et7Cqm4tM
mh/ofISM7sS+vxdHtmj4x1BdPlb8b9l0Wg4xvey8aLCYKEtIsdiHnr4BfTTW7mg6
gQD6kpyl9a2F0YWa/6pwChVOOtx1LPQi7yxJ5JnJR6TmBXecWGhpH+a/aKAxv3al
Ho04gqMPjxSsJpua+zN3VZNfjTVkfjV3MboW+f5JFW0UUhkJSbxpOfmcs6LYicYb
6wKIgigCE+7/y/mqHvvaORL3kv/3AwqXW2Xy7rtLcT+OxsCxVI9Nr97EQvD1KJ+B
slH2p3LdZ1r+ymedPrFUqcNuqroUBcDWOpZnFvxh9RRYVKAjVQvpJYRzlrGiQKDL
BG2t1iRuwxTF84HFvdINzavtvJFhDeYl2d1Xn3dR10zxb96vDgiYYDrgAiZPbzIQ
BroZM/rT++/N2nomBPi0e3B57sCcHPSRnDujX2ilHFKCLED6dgFFDrJjk0vNFCpK
qatZNLAlNNrYX0HxWWM/nDHOhVuA5R7J9/WZHjbohZkU0JAXKn063yq3kbe8edwM
sqB0MNsHcx0kTkEF7DM+Vu2ebMa77iAs6uv/HwpLI0Ooi6ZQOPXo4ehB0QcaZoUV
nceS2D4Ak0dsh1Xt6zvi0F8d2nP07h6HiZ8ufUNiw6mB4mhcbMA0lmPLfgn/i52r
SrUftYArP+60ypTVx9l1fZ3H9FBNaBNKf9/6hVjoR37t5jIk/yAjZL7/0f+yy5V0
LO+Evt9AVgkga57x8UhKq7znKXzMYsQFW1Ha5TTwqr+Ts6B2+B53bKfqN3VambNE
F+PmOwvJ7TB2CokekNBzqNFvWcgFoduA6kC6DFGAVQdipJ7DPei5/3dwE3KW+DuK
gso5GSPsIkKgG+CTHXjCBfPIrKnZnEVIgqq8UDTE2l+zuogeAyFH7Fs15btsS+/u
dnA3EA+ygpwFoN4i0yiPOVjFgzcRVBaUEvD/GJBAN7PZCdALqmt4BKwcGimJS0ZO
7augp29QjCJ+bANZzHXQ6sGkB4iXs3NuIJC0mjEd6dDX52KNg9MikqjnlAGXCm3I
6jwaRUWHo8I0ho0K36qB/xQst5aD7gMP7NADyYuTj3Ug9/JWr2qTIn9KERgAL/hF
jX5kFjYGs8j/SqnbyOi00Fxb1OJxlBZz/juYfdYFY6CmLREj8m6fsoJqkwfc17Qp
E6SkkGRIuu2YrIMBCpI4Ij1UUf7gHDVxMB8C4n508HENNuMrAVTnt9lRXVeo7HUS
sQVkb/Y6Ely4JDlVXIGpde8cf1ptfW1OyZHkLD2n5TDxhiqROWeebyUgc1wck6eI
4l1MxTbiTmReHE52SlrAutGH376cemG3/KXLvEDJKWR2JKXmX0mJWdDgPwYpPArm
+2elhNvvNog9tJ6FD4xIwA/WtWTcC3DKsGhfPsgwfd/Tlyx7OjAl2h/dkBooTT93
hjMoAnFk2WJ19MxKaFmSYdQIWjWCDvgsUt4rg6GPHxzOq5S8k7wm972tsk3MFXd/
UItaG1vbUgWje6U58Rvs3sWuek9K29bDdcZ3vB8E+j1qiSxbzgMtpe06htKvbKRl
elI28ONZIJ1CPqae1ElDrXk8hqRsWTnWbX1o9TsY3N6qHJB9PxFuy7qGzkOhOJvA
O4/1DOWqM7H7J/VbwXGHkVnBxvdDkkZaeNS3U6SIBc1ePfkFluKQS+mw0iJ+Jqur
7zUz5yd1DzycLSRXofxQJTvNuWDNcz/CquBYo+NHeEzjCyNn7Tj9bC+IBoDu1V05
pIrSNyf+/G+UzUrVb7osvnDfvLfSjKdG6gq+N6u/dyGD18jJpGxJE9As5ctXS15b
XUxJCMmluuWfurDhlh4AsU+7y8DG93u0kgIRTIeMCSVZHdLh4OSHV2JXYb0Xg3Dc
GcEZ7+ZN68SH8cqggJSOrkRefVSsypx5DHNTjGR0S43jYhLyzyE1dWHoyfJj/bv2
OgTAUMAVRiSUo9PsGGdCLHPgRrZGOZJbjB0XoNoAIRMAFtAbbHh0uQbbIggbwNyv
/SxEvycLBpSAJXYfPlYepoJPwAax9o2uifKqD34w4Uq/3/W3CDzIqkUynmhzhthZ
kr/Y5Y2/JfmscAOvAz76nQE1xf7jabXn/f7UXBxscazrFLL4BNXaD/nboKJ9zs8V
ogtgumhhQ9p7MgA7TZ9NZ60E36puQFxATr4+BRJ0lGMwUM9kekA4nmn/91pxwfTl
dRzu7gWhJ8qiP16wOs3Xdta8zyyy5qOl/x3r+xtKoB6Bc7muBo24jwe+fad+sgNq
u3C7EGeaqcxnePMNhfPGk6ym0if33VtJUTEQoM9RzUUIG7YG949/4Hf5VSGvIKZX
g1bCTG30aV/i0n5DK9jRXr4B3aAvELaC1OFKmDIOtZY+YKaX9Z3zsiuVIRmEhdi3
U79HjCoxxC85p45rWmKjy8/F131JjHflvtBWBGPl4JOYPkwbiqVelhBhU00Rk5/0
5c5q41wAlphXH6CZf20j3wAXatT1eOY+togxFDo0P1Gts1aRaqMqI6AmBvLreCOD
W58ZyvGizWlknGX5zJAd3iSeZroN2K4sTnu3GARu16+DHD7Vp7kSzKfpWKCZcDoM
oArUGnaZhY7a+nVOb0PYc+RCUQhcMluomV69H2ybZf65gEkuD0OVTAG0kvfKviT+
1mYtiL308cB6P/T0PgkrD/ULU1CgiiDDys5xfdKPHc+ccoYOQj17dtbgNqQJTyeW
yRgd788U+FVyaQY+EMrdW80Cp2mSWdplf5I2farsexOngBaEXcOVlMIa31Na1kz3
g+R0aMYKzOAX28TBCdwd8erRRv8wxvrr52sDpbkAHT6tKfp1C9Uv26GN9wjJrAK2
Opp/kX/EDgfqrC195B5J2kVQJIH2zUhprsp8Grp+28kHBZJCOUgn/6WV7bIPIa0s
IfEkXBJwA7zyJxyX09pixudW4bK5OizmYeJ8ojEYHG+cOzdz9cD9CFXUe1esa6UY
ZQ/jbn5bfZbT5vpAB/yqpGwDdu655ZUBvCMxlhKVXPuF6djdCuRGqloRzFM2KV8O
fQ2pu9whqMJTdrOvq4hcru2kcDg6LsWvv//g2ZyAow6i2mEdbsY22Hm+V/n4KVyq
r3tmBNJBWz0CWDO0EkfeWVxmuJc1QkElxOb3MHlp1enzoILchTnxSu9KPwRS5i4H
BhIMhGHVuszPgnu28vxABMFsr/y0eGMtd+rG0XlM+gIHpGH9usl5Rilp1LseD3+v
v/300Q0aLJY9W5lxO0jUT4BfW+nXc8CR2qjwJj65KvH4He89X4MZy8U84xR4Exhb
rnEhqYu+jng+pX9oG4G5a+0nnYdW5hu2ivfRKjckxF7OfHOpbbZbUWebgwvw3bZN
YFNp7OuVcxS8yNiXZfD+vUD9kfRDD0LAbNcMDUVtgxj3jbB7k9e1hm4/9ms/3vW0
esyxkLADMWPhGzm15N56+Hef8PNFwbGBJ2OjqEd2awkCcqDOi+QInQBpwNLhzF2G
LAYrB5qDMo/qQpJHEEZCV9BX7exG/VWWIim0b5JOzcFj0YYa5mDNZlB6tenvJGzS
CE0X7WU1r6qjoWDfUAkYPvbUI+WcRxz6aS4BshkZed2pkw34nAOt2w20DZElddo6
7A3FfKlmPeynhsSj2HTivQhCGrS4lGR1eUZczPDnRceKdvrCiIh3GWBSAihyGaVd
QHNxKX1Nb0DyOnOMblQJVi3N2L3jAdmG9M9bgtGkQ11hkjIDM6n8TO8PIq0ksdJc
3Dgx7SQS3Hxao6SDsUtAaFkQiWA95xi/7mpqJ8K00zxLqU6nBW92zvhdz8z0kekd
AMryfnzxh7GrsW8pPBRLU6rvGYzxVcqq/C2pxdlLtbmYX8OdYRPjWL9y9m1YNWuQ
sGgzcN4w6VuLo3wyCPoh15QsPGzkhsNIMdrmNmy/T8Jb49j5rTvo78ng9ha0ueAv
VeE3RMO3JQrhVHmm2YZD9wLmDnMeiqStp3wMKp11FW8NoU5sEf5njmsM6wyTxTbB
g3tjdmJuBwYK8phuj/+B5t1gOLZOlLcvgvvHQk5nLA2HT/GgcM5usY+P4Tz9pWpR
Gx53Yy7cL2QLXJgBztDvVaF/AlSi7mH6zJ0bAq5FqiJrxoxYllbhBVIkzGmFlJt4
Wqhw16RJudTcBRWGdpYeX7awubkzN6pGANIG8f0VrEDePsE+9qMXijAPagJY/5Ob
0Fem3PmU9qWJ1UvK4/yzjxxkWGYmPgIQxP1Ii6otJDiKHRWzpK+JCseOUMTWRIuj

--pragma protect end_data_block
--pragma protect digest_block
HZI86am9lJltmqH0J4ESvmlwpwk=
--pragma protect end_digest_block
--pragma protect end_protected
