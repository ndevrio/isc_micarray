// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
cdOSoiheTGg3l9jHDoM5LpNNcDckFNessWWLrnbduRoL4HjnqqwbIlE15vkIp0PjDNO6MZV1l9Xz
Nw+XiiBIcW9/QF91sR0pxX+cLtnHWQ3XhwMzNWPQsr4NU+DNobD25IytuY8GTx9G/8jsH4iA9/Na
CkoP4+Wv/z0WWgkuYzDheIIEakZsBIfWFQG1fz959/zRGmHG4rIYx942W84Bk5sYTpgzMw7L5exn
SG6DSQ0b95JKI9BU9agFS242/ABe8cnioHRADQP4ORZfheh7Ut+1ZEaXXdmvXIz5QutbRf0O17a3
j4ivQN6ymN9YXK77vYhdSL9ajXfuZPcJuilyfQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 16704)
mmbdG0GUp373H/rFNcWtndo0asf+JiidJSufSt7j/9x8DSkkj1cuYObMUZpQECBtkqm+BOPHAdJW
/JxbciJR7gsZp9KoOPaSHbIkMOgNLCWQVFxn0h4YDZ9W9kgvQUXhhVM2SlMqxwxqwWnqLpZy2ZvY
oKH+R/SJ3HT5IL5LGO0c+3LxUUVsiRYqLUBd9W/KQfzPTgf92rgPtRzxU+vZKSI3Rf0C+Sx02bGz
Dit1IAG3uYOZsBHu7SgTb3trBN2WuUXUSfcLY2O88XaH7TKIQ/fsDP7ClBOFD79Qfa1aGyv7vQbL
o9nlikGsbbu1xPszclt5c8bow/ksli6EFWUI85lUeSlWglVoBBV+skf9tdaCzLHGzHxMv/h0kWcX
clHCq3cAS6DWk5QSPNZ8kBzJbCH5MkXoNzxjvnMfIentcSVLb0ti0WCv6CbFaIx7qIvFkRa6yO+Y
idXyskz2lkY4ZMY7c6vUAnyR1kJaulJ3/kodfqR7kyjBhAwU36F8amCqDYe4f85zgsP+8RsabsOh
Wy2cdwh4IfOm3I+ef987P/i6awCVpvHion/XhRzrLKGCN7YcZvV76kpzHrrWv/H9/iElVdn9OMT2
lxo6IRtMOfbUqR8qHy/H+SLOroasIuxf34kxYFnwYxrZvI3mHzVKIImQD0iJcHC8n52FaEUaWrgc
lZMd1jwZLDM60/VL8GVhSE2bpCR1rly8fI4Gp3KZKEVYJbtnMkqBBsUvkPAwgUYbhs2IXBCqlkyU
G6xqNNUUsFgt9TAR8SSjvXtgUW90H6BnILzIhQcbT0/21ibYgUpgx7O3LVgAljFcHLj4dcNUBhCr
F787nOkXHKAiiPULpH2OuIMHwlwNBJd2znDU410DC/mFf0RCRRaoS/MGqnfvlirk3y/yKpHN2ZnI
YDfi6oHU+NR0HA6aLPN5PzafFbA+LWSUgkZssEY0qHLA9VaA+YvFCEfUvt3JlqLW4csss4Mw2xUk
Qr+FqyJmZXerdUBHYwXsOhzoe60eZIkbyvLRLdp43JftUsO9/VGwtfUdo3a2M7qNhRCL/yZv+i18
40WfFDFodCfwwJLTovR0muSFVgLpMeoDj48IJOvg7SBjlRr0jb/mXIsQeNKB+hp/IIwy8hCbVHr0
ZP2bRF6MdaUQTR6CLjB5908VAmSghnksS50XU+RFsKoeBAV5Lm+DChMUauZw0oMXuF1GK2qCicy8
GCHZBmTgBLg/U+FIWGOS1pnHPGrTOCC1vY+hbTsM/TwPxeOq8fGgCU6BvcuH65JB6SYV3eS/kAnT
pm+3i0kMxuuiRtV5i7U0ryh5WjvFCq2AYns2awI95axRo2Tq8RhbuUrmntYSB6DBItTqc1wUmOcn
lPH62lymH4yzF5IPDycSYI30rt4uCb4AXTe5vjyyhzAkS/PLZLz6f81oqeIuSOjO4rwHdgBs2z4U
Ii271gCDKqsD76zQ1nwAsgRBbSa0d5y8d7ARyE3/eYK0QVSQ/eQBw+1Ftt7SLJHKiR+TYdCjgKLz
PYxl661kuHFGjChBlyexnEPvtw20mB3JRsV4Bh51GAd4dEa8tEBYMZBY/mbmT5KEr8S00jaVP74B
GrSWiWgFpK7LgMuav74bqeMRD+Gyxw5V9F/o320Khgyrv9f4LyjPEpHQtqvoN9114aBGSDOfHP/u
Gquuy1pwcVsamAKzwYdQC7FyQ2AcMBdb/UAnsdc9Ml23WXA2kks6xYhnO/pmeVn5dwcsrEVvjNYP
Az+aehl9u4RFaih7MdwL6H+lwSxPHGZRBfFUtgl4agkpNd8HkE05fqdvX9AnkJrTlEp7IwvKvs7a
ZROa9ElWQdCNTlCnr6uOoY6O+Xc5X9TTR2yOgZW+n/sAarYlahY0xRt4cTaS5X29vjSZbyC2493s
ROdqVD0AT+0B4YKJLNY1Spaoi73mZzxlI3TuPsMzei3Xuq4bXQ6ZER0f06gKqkNR0RhZeYK8Tcre
SSun5Ooinv/eUx9DbBwCmSzsJwaIixD5zFxraXwzu1guUuvZrR0Fhh9IAkwiUsvSfu5qfE48GGoS
dFAdSBAK1Tfo8QNHMPr7jOtM6J5DRmqM6VJ2EzF5nMTqO22SnfQrVuZWYGwUdiyZEEW6BICIqutO
UXv5aiVeUIqeSUBamdoheUXbklBl3U0c+dI+uxt8vgFRpIAfImiXz+kJXRzHI7EMAR2DZJ8XMouy
vgvGFJsbUIP+HsqObrVbyYqWcGTplHPF+flh35UnVtdMfkFHFcC3IlpvKurPxmHzUYjdGJ7Wl00D
Bk6osXuY+A8La9dX213I2Tnf1LnZE9ou43hCMfkoZq2zPYmWQqZuQTWi+lNKigpmYb/HBP4IWnqM
AiZXSuxRo1J2ssT2iEWGX/YJ7xbe0TKChttSPVPfkLt17LGCl0j8m83dASPckpvm003f+VO40OkQ
rIzjNo41fMWLe2pjyilpH5z+7zE5YcLBI7wkQMzdi6l/Wo2/STcvyXBavBgn5484W85Wn2zndwQQ
bvBuO/7Ogh0ZqtdZOjdr6bszi6lBpWjt246TT10M75IvZeKn0ZzXSf6E9HKwy20Mcv+YoiUjel8Y
4SuDRQC+jili1T5NbWqtLBpRSsT8++03Y4/lym7T9eey8kHsr/71uhkm5ZKXv+G0/ddbCAyYckZp
gFKyEnt11HX+4dJnqD+KZxkohTNgKvT+c1CarUmvTQ+cyT0x7oXsvL2OlQbvfk0zC8mqGPOmd+IR
hKmDZn+Ha9dKyBSDh8kEQ8WnuC/I2b6/FBDX0kYxF5OQDb52VIZLFyRvJDCkSScPACgJAqqa+mJA
ICc2xTUts/skwZiWSQ1XpvtPMKIfa6sCNvTjJW7544qwRY3yDlwAO2xoOU6EFwMPI09/SW4PJXeM
uGkL/MwsUs6tIudgDedZbAe2YrBvX2vMccT0yJeWH3783JhqYR+zDWacJeuydCXB2eG/DyRYlbcp
JhlJ+KL1RPaRNWtg8hkVYSyAjTSa27Wf9WR4DH7lb3/WT4mrTPVH7QunobhRyjfOKjczKP6jDYnb
N/caGPRvhRm8MTyzYrBooLvazzIqA6q885ZgZifzG2/8a3OMnLDTYHvPoDfNucY2QEjTMo68b3TN
zmxaXfmpGmg3nkvgEVUOew0udLYscjo8JunCtPIzuqjcAoXnyhslbcAJzhA5Ma55oAd1kNzJp3j0
vTO0WrR75XAYzyhP9GPyHdpWkwJVZPZVt88NbzshYxi5flY2LpiCHyzj1+ZJErJOITPzIsCrxBNI
KvXd6NDvIsDLTc0aYfIHg5tAwMYscIdocA0RZRlt+NEWy01MR30KLe2YSiTxNrrQb9k5hIrQ8ts/
wMrjQgNph74RnDa0Y42wkYGzKwTgYuTI3FgZgMFGt+PNvkZ+o48T2b1o0992xkYauEY6MclH6haG
o2iwYcrnr/DjdowoaoMhTek/vnggpX97fORGy2QfTbG5g4MpYmyP64/4/Arzozy/ERMEbYq2NqUM
CfnckcHuAg48E4p6uXSe1HsYiLXMwbHMrXemqMQu8n2gQdr/FnRqHKIOukZCrjuihd2IDJH4gWAW
/80WyQO9l1jwNI1a8V9ZZHuwaPQbI3hg9MdiYXMY8nw9aD+PcuirXScXpH00g9Yuk8yu32XUbPlc
1tgAEA1dajn1HKMBpnP3tbuyTMsfEkKErf5M3qwUkjcVNdu8BvENJWVjQCkExcSvD92UPSX4vLWv
kVKsnPFhOlCjxvM/C2QDnlpjGigpH+v/NWr29PmTQebPq76HpGeelHDznnPwOIHNDsGmg27hKWW+
O0VC0a//QP7F1BphijDWn+kiw99vuCCmbmi/fUcU+7B/jk9dLONMx4yL598jX6wbsVYH5Yteds7Z
1aWOiBxcxDaHUM1W/6MT2uzUzoZP8pxnZKpG6MFBn0Iz67eLZU8WFj78Y1MUFcATS04xxsj1ReOf
GRzgbOqD64dZI2opeC1WZ19OVre8I7XNgZ1KKtFrLT3nNc5i10l2xUcN1PTXx8+5ZWE5kI38Rkhn
QToMRrt5HVE7mCSD6C7qVVUM6/RBoleofDYs9TWIwKCBfLovhNxSmz9JjOTT+KO7wgH2X3nFCV1H
2ACW/+Ksb0wiElU+ar2jnDiZE542+2KuY7HO2C7GUNIUctLcjnmeoQU2N6BJaQga+1ap3oFkQjiE
iFG5De0rPfakKDjusWbxtmrl7592X9fwxoxDS+E6QJbY/w25JOFjNTWwlbreuisJsq+EpMGjgE4d
qVVtnJ2LRuhNHXSR6bb24zsFC5MB/9oFpzQYvSJGcZ86VICFrpKBhZpxmpltFRNyyu78hr/vNj/5
Hh97UgFgH/XVK1UfrDa4t6Ck5OeNiQy0oZh5rDJyvhJMJg0ljTmyB2niFpmaio6j8Q5WFkMyHlvT
94DU5WZ+bABxkEZNXWUx3jIuQCFY74zufXKvBZd8xLtXXacOIA07egSFpst1lbkHlpU46NWWVJW+
tS96/1rChPiwOe6a3EPJ80N9bWi8Cs9hD0AxkvLL0G1RmraHn857xzThneW477h49KIpIspGC1nn
lpGdRv1h583QyjVYUOMuB50trMRIju9eW0w09H/ySMX4LltrXi9TQw1BRQzfJlaYwupcJNBq4miA
FiN+3AAkyBkHlBYfY42g1nQIMJx+EYkaQRcZUQ20DPbcvHFpmAT4m0mOpZiJyd/80+5wQTF39X6B
WR4dLXzcraI2CgW7Y05NjYAks+2mRoQqC2Axhd8wW4qkjXMle1To/ZJbHJuDIFSyTiBvEC962vv9
fKbisVyFAX4A1UUEH1KKqV70GNnQC5WBeQKEif1IsLwdAoR7mVQNnd/9i+bapQSTKjdDdNkdQ8Qg
g1VphJz+AXiIrAcAiQI07VsOMAsSGUxOmw2Hom5CGqM2EMkARFipX1S77pMz1M0LufK0/fSxuQkr
LY0/uzUpCe2Qiw16znG+OwUkJ9uYdOpXyLZOhkKxVivO92Ny/St5PNZ3HRpTBtHuz5L6U2DyQVU1
lOSUaZICedGX75rtuMgMl58kE7+Mifv/MfSuihExS84zo/hmLGNXmclb8UjlPqhpa/2x6xV6GPuh
0Nfa3LMU+cVoCmHzEiZaqbOcz1fDrcmfQ8YNk5VBG7qiLyZfrJmUlo2XkmUEYXbP4MR72dEj5DPG
wlMTzdr9EHuDrnetV9DS4bLZJzPBb9cmlYYC2z5CqjH6EeP3xFeWKf/UvQNmZZq1mokiGhuWEkbG
uFLjJ9HePKVxX9i62FPwkls09EFaX8RU1gyIrkpekxnWmH7rwPs+wqtKsbovQmY8+Tc+TGE7R7Np
XLp03zgEt6bkGR2dTxN4xHjdZTvtAs3qAZbZXZRAb8RgCgooeSVUBhClGDpgbmikJ9CO5+QrVPZz
IKiBMIpBb2iMr/u6ws5fiTz9Z3Iv0LGdOXMsZW/Ku7doW1dAsOSiRxZydNdzB41j6dz2wExoSMKv
NofFpkyMC+87adb8cee7OQbn3sXGrBWPLqjT8dBDVd+c91yoHrRz8DiTxIV3eP5uDVwZx3ii4TP7
Hg+XT4GVTSjKTXaWjvtrX/bEv523rEJkTd1HU90yEyNxzk34xGeGePaLSck8BoCZf6VLsl3FWezP
o7OfpEfLLpf42pN/5IAObaBZcP5DYto6pbYLuphbYx10+jy8uqehXHSOWwp+g+6pAzdY9aBIjPOl
bf4AJNSnX/NPLxSi0kvJIEoLAMbVJCYuulezFlJTGTcxs/Ek/fo4IjTAYmoOg+OmO5qcEyxJc+8Y
xK/cTdf9/b3McUGiClUfUueoDkbd3zwhLopCLw/Fr3NsQOOW+7dcwUkHJsr3iRbBGxsIcordRjHF
uDI1NfI1YNQ/tsapzNEp9H5j/NXn2gM9UMtFokf0xmBD/SQXLLaEDiewVmCW0jIQeJOfrMibT6Qq
3kgU+q/wsZbRSWjVfYYXgJ0b5T9zSbMSuaoxXu2TYENYq+aiAz+QkS53NIAdg3daciYR/TdpZxdv
Hf3Pn0lIdTxa/vhSFaJcFdEPd4saDuNb9smT6EPY1gPZ6Dc5iffbIOT9Ant2q5Jy4KVwwVu+PoMu
u/vVFD/RmU6xVIx3UmH1ikOCF7jk5J8HQjI+lm9IowjA+Tsj2jTyyGVN0Ju1N8anwswpd6wa/zlt
q91X1w5sgi4VLevfYmmB42BRa5lMEaso0zlEifTIqNcDZUwiEm+7LAHKt0Q/b3J65ldUMvZI3DAH
JRuaRZlfJb6mohQRT0GFxd/YqpmpNcDs0ZrX9t+1bKB4QpFouotsEL5hFe9L1vvmAgiYT75+2Gpc
s4ggoJP70oQQyG6rz9hdXlwGDhOga/SZGwGtMix4zRrk2mInoRqxup6zqPGdHr0Htc5kWER5ocoo
MxJMbGXUIijOonu8IlpSZwCliDWJLnmv5uHSme0CrcF9jLijwdCUrIuPkJazjJhEFwduugcTztxO
0GDhd2StbVmeITMFv/2ncGdIp1dlm4NShx3uJRuR3aGWSRksr9+Dj7wxUWwqXFiJH5i3ESzizIE8
oWDGVTgqKO9YFUbICFtTX0xXSHniEplhuk9kuiP1g+cbZ+JKInzOd16E5ld4HZpS0c7qlWKpPEVM
WAg/e0Z+ZqOWcXntZ54/6aD2mRsobarn7Lde/8FMiS+vnOE2dyVuYktFr9Wp/NSWeHjfyk5q3QO6
MhYAZJYP66LQMFQa/6RZqwVxgSYJyAvTol1fREYAhOJ2r730bFoffpfG2uDrek+LrJAuDA/qYfnW
8wYoDn6G2dMX8ylbzS7/nEmhdUsRTdsyxevQbw09hJdo4vIcYgLnlRlVX43i2QQQ4xNvF6zM2DdK
jobOq1Z0oKjm8EgjpdW1Zlvlih5kD8v2T/AUTWpZbqv3Hbt2FXEZc6URKDFJHC+91xSFw9Q4x5Ht
XyM8CZniRm0pl8WJLm4V90gLRdd0CZzwXfbiWJecXHLs1zESjKmuazISghH+6ltKMEKT747krE9J
A2N6bsGHJSZCimnJz5fmY7A9/Zxf/j9jnOWsnmbCWPXQX138AwJRGeTFmOe3Zebw4OdWcEF2BnIL
1KO9tgJuAXV77EWzcvcCohlqm7pGWusD8HasoxAl9qXnDTwIjYrUxJBgbQFNl0VwNoSe0+7JLvJc
vwflDGwXfz9yfC50IIxeQ8Jq0GrXZ6C/+9yZoeH67N9ulFvUKgJTL6IxBOXv1tsjmvxa4c/z9mPh
836CJ9CADm9cnju1ryVIegTIjV/h5w/KhCqyOQcvLDq+QTNXAiZFqW3ChND2DLu/HlBtgwoS4/tc
w3l9L0GZjtGtZvQVP/RyNpk9yGLoXCZfVtySt/QNoXljYkF5jhK8GY/0i/VTPFNeSmtKWcuNr+dU
5TJUkBxtHLL7j8FY2oD0RDwV6VSx1sgdM1PnewxpkKKzd1cdc09Rvab+9nij3o9R+1NGI5DHHt12
T8jDIIQn/jtfqS4SaXhtXKqUNpkC+HZZOtKrw3UAcHl2Xmw7Ds7nlwON0vFoWyYEqNj4WHDnD56C
yRi04CagqB4DstnYzcPJbdAIIAmfa0Q5FnCa7z6OpSdJK0Eo4EjFTLTOYslmAK4DQ5WgLXbIyWbg
nTJIHC6DX1YoSzKhI4iM+SwTihny+JRJZchTvow+02ANvQ/GKWGVAxH6cLejl2uVLhrbUTKb3m5r
xNKAgXqVf3u1ZBdHz9nSeKV3GA+KvK+j+M/NymFbPFyLiRh176dtFtgXPlrPk5zaaiB6uSHkA1O3
POJWqYS1foV6D6PiI1MUjv9OG62uLNuYHu2WcrgMi82csrEnXpTWL1rdug8le2PE0j/MNB2QOueX
Bp54DEBQA924K3c9jJC4mHsWgjVNT7cgF3t9+1AJyd1JaYLlPUoyWQcE2Tc1JPTlW7vHSi9j7Pra
YtJXG/Xv0/G8aNCYqqsWKJK+fY7ZC9KQwYF7eNV97927VZNk+6UBcFBxZ73YbQB9iWsn8kow8mcS
ozyv1X9XuYTcxoygbZlxZ/mJtnUreOWXOYIR4EgkY2y3PC7AFHTUFLD3rt8C1P57Sq1I1C/w9uZw
jNOCtSKKyVipxsilND9MSS5UPwY2OuHOnPGaF+gpyVuMECF/tnNCiF3Us+cQ+5zDT/3jfV0FzSLT
jdPltbvUXcw2I1e755VJm2C1HPzpgmkPWJeqpjsj6CQwz21FbBFbq7pQ7i5yD3wibu9FgRsUPaAL
Q3EnwecnBw538csotxmLGN5/546iaqcNlrVAGIR+hX86vwVeBw8xphbXVWNUeRWBbCv208xTBXmf
t/Gew17OaSn5A7uqMhkTfctU6Pr/x740vTwjiXkNB7m1cIfwIeg0z7Blja8DxyUl1IqTBiodccCO
ujmeHn+57xjWEuaJtJ4KmSHxcjrrmujoW4JfDhGjhPtxBfXbbSzPY9moE+o8RGly3cEy/+ifG7FI
i/cko0vs77dmQqVfumN07gep29LK7yQrC2H8Ev5p2LbFWyjcDBj/LrRDokyExw5/HYFr8UhPxWTq
AKKO/zPl2729Zt/y+GZ80Io2+MsdXKxvmoDW427078udmYI/4Wz6OoNS3SnAUijZwR/XxdjtBOR6
Tf6+O5RWSMBP5Ob4J1JL1vcA169tsccK06UkNOTU41BAS9/ir60tGAOvd4VLanbNp0gFGJshPBAX
9QvH6dGA9h6FUhuiiR4jwvkGT8bm0u7hKC/JsOoLad0V74cEDgLrYtAjLaji9olQTJz7h7DURCjy
LCL9/IvcZ7/rQgPCM/D2bzBJPO8/xYtPmWj/nbq8C/1y6yJ2JNRO/o6Cl+SXkM+/TiaoPDVmGspu
zcIy3gL1+MUniMT6ZKhLAZMc0n4j6M4PdRCdBlipi2gn1zrNTx/65fyeWW3WQGEvsb3CZbCGoOMr
D6nd9in5q+nCI3GmRzSGK+tzFW+CkjyEAKYx1VMMvQCN92u3lP/5bmEeNaRTIZpTJ2d6k022YlY+
hSIboyB74lERmHsw090OmNlLFHWYR+XmQlTJ5l7L23o5z88M4x6j3DEdv5xv1RCEQE2sdTHAwMbB
z3sltDGJ9Ud9OCNweHqxjLrDDGaxNaIqK/jmhymeKQ2G5TK+n4xs2z3hdQTvMLqwlo2f/uxX1hMp
jPuR/c0myAI5nPzWJV8l7ibTHFa4seRBh7Bf8XDdSfZH2I1h7wXLyiPG39C023qaQSIhfUMOWeEK
Jwkti+L8co/t0GKqga3CRDQjCVZbe8Tz9cR+On7U8lPrTiVUqtWToNY0nBFqxrWWPp6ymddeVjiH
VfM+81o5ydPfSbEi6zmC1OhGSqYaEDrGzEkaDw07GVRvHQBl4y42x2mUqjEpE9BWarjUFUw+74ZT
YmjWau4tWofveVe4IiDuPAYUBPlQF6RVbyM+ns5BGCls+mVVxisyhFjL7TgWmKzkacP6uEJN387e
Ei2Pr5ouZfxxlQNsw3/SpQ8dP5aFadZCemWS4tUduEW3dyuZ0Mv0Vx+iZ6CwMxGCNG/rRT0i4A4x
s/j36Hm5o6J/Xfk/MT8y2fWHZKY0gZXERnLbH5Qd8pXtwdyC8q9F9rvUQ9PR6PltywY20Bf5uGo2
8zlQr1c9QfFoN/SrrKKmQer7EdhlIJuT7VnY0NZh+fuQkgHqnvWo+d9Tyet9zbuJotEeyq+2Gq2U
u0k2/JIT8taXQARyaLpAR/ZAWmqA3LHynO+20d5Bv5oc2sV/zZznmJ19zHjKoIMZKqnYkjIMr0Kr
JF1U5pyuoreCUiVsI8jsRoYJSg/z9XJNYsaE851oxtQ7L63LztUK+Z1yjOM/8w3uCj/VuSCFucu8
eF7cDB8HINIDvUpElS07g/HpFjqw7C3exk9tYDfMt7MYuDrA9ULB1znqwynswOhRlqGxtvjLo33A
7utflfkPDTWu2BmVnBh47Q8MCNHT/2zOQM4EyXZDXaCxAjn9DCrdbIHPVLqTKikvJsr8yYHWCWpG
wGiZ6Nq5ZmNcXlmmKqEEHir4Vvd4WG0xE2MfDoZkAsyZaq8P+KHgomSOvhLDuJsF+HEeotqF8Gpi
jEtpR46ui2aqogfLSsxPczle40UMk0QerFGNzonOaKv7M2TL9QwvDpW95CQrLcgOBzu4QGQl3W/1
zV88IbpTcfXU+q6kdBd4wWaskdPBd2w2qrB+hPLyK3lavWDk8FXTI+dCtIZqGung6Eg8NdMBLKeN
ew8BIyicgG9scSK5l6bDcDuNt63UV2emJ0nCQThQ+rTTtF4+qmvd0p4kgnAd88qCm6fyCUqwAd6A
g6FNRZbmEvFJj3FI7TuxTa1Rq8bgG1ZEVoBx9aE2Y/ZATGAzsLx4fMAtjTo2UhzON1KlwzX1L+z1
7PuZKhJedvWBfWE8zEEcFisuQIIV4My81yZAHzj67Z3wLrpf5BLZ5S4JFNsjGpozQe+PpZSOlGqg
XvGD9AM89QSTVwEdLfNIqv/E9A+rQ+/qVj2xV8m92ojspem8THohsBR1BoPAmRhmkvgoNawOeq5O
7kOVi+XRV5D7EivwSDmazM1xOabTxks/943poJbkHdom3YE7BEiJPJMpxe7sI4n2h81VKcBOIJta
3k3YPQM4inZtPbROQeMICmnXkie3MLkWj/Fi1J9GUCjIEhE1FPatQPM3EFYeLZDZKQMP0/sr+eLQ
aSftMjFm+Uy7f70XyhrtFsq/vzF4oLoYiTA2Xhwj0TSnWwp75zqR2o6o4U8NXLrEry6nqKRd/NgV
8C5jYkpbe6ba3KH06to8S57D3sZHw1Qx3FFfBm9Cl8lAX93E0ZuBiF1L1oRO7Pr1xXZflwS921Ju
6jPLV8NZFaYzyjdTm0vyBPo/W4HUEheAxsEurbaKeUHgyRRFbxXkZe43WT3gpNFY6ISBGp64f6f3
U3lPomYCiwS52JVs4uGBCCXIE6H9kHgairztbALFRnDf1EgMIE1v0sPdvNIjdZG1dBVuUUFZhLVN
yYAId80wPDmbld979iwUlRU5OiRzZ6jfzPTmqlhiDoLsteIhbcW3gSAA0HbnF9vGJMCkrBCS2nlM
AW3cJvq2B9V0Sa7euLQUSSfl74IO9rR8zlNy/0CNHHKG+VZWbvKQSeF1ZI1UgN/ta4HnGAW6dtos
UfRhXtkXV+fYTgCfUemJIpHb+hvVHuqB4QYBMdm0kMgdiVHgLKqDiwLH+Oycebnpyz4vPPrFRC4H
Y573NgNcybU8lUcK2QRW9/+BGhz9RBs28ScFnqrv+NQo95LQ34nLYtfFA7qjCUJUwFAGDBcxwXuz
0pULhH53CUfXjsS7Jvsm9ScbxabgXZrLMThI2J/cnX+inDGJcXg50I03FirXbn8tMyXC8XOQGaTz
3l5TnAlo9i+kEezvO/kWU9zJiFFoNybkFoPPZGa4S81aOOndnbWemohLziWSBLg3K2FejC9i7eUO
5ItjPsrzWvVMS/gbV6SQBkO+TAU/tg64LsMlbVq3pqRNH5r7avO0sa1zCwHldravAR1/BEttB2Cp
etzF7GQU2UDwWm9NGpjFiZoOj6CKUTncoxhmFxbdPqImMxP9p9owzXTNPHtY86Mlaqec/rXnUgH7
Asizk1OPNXpA+rZQ+BAMjZfaKOvpGxMOo90S5Cx9oifcyIM3ra2bxxmCOn2wphzdyrPbVHaTXlWZ
JPtGmpREvWQKoApMg12kAQYeLzbaLRpDmMheqgHv5r/48E2CmMZgkJj2sphJMFEfz/CO4OLcISQk
pHQrelhJNrOiB+GimJ/uIGwbZ172Zu399sQvmBtMY/5liRUkbhy6BjC3urSEYUuTdc4/e4uZdmkI
9uS72js6xnahf8W7/0T6V0UKlJ3BvSoZj/aQh55cjd5+a1z/aY28ne2aCw414CFvd5WEUtqMKUWJ
BsbttaRRa5eorgO0ryUKG+oWDEKiHj68QH7347hAk0GhN4+lB+312V4VzFpR0v/ynYYCm2YdwC2n
SoUtz3IHyrVMHiozjS0sEq5EydJ+7OWxMWBsWdXsKxKzBzXaPntGntaqus+Uunsh1EF8uH/9j16l
A756+9vqytg3u8YLw7TNUmJSKA133hR625OU0R8O6E/gBuNiVjBba5CseOy6Pkz0IiSyfChuJYE2
wtqhufthBK0Rd80edhwwXDU0KAiwcaV6y+GyDSi8U8w+wwGe2oFUqE0dV09wtFiDT5IOmh/J3niG
4U3PFRMzp9KU9eVbiTEvukWLJKQPrTMLRVxnd6mwY/L/Pm0G8IIHm02GRkf22aZPSuveqIqzUT5y
ZzhJAqVmXcDTPzqwkIJj2N1klvNfq5QLcbK4SFpy8x0Hc6KXAy53le0RwE4u6CChs0LHNcjxk3sO
H6MY6PiYpDKkJVdVgytw7Lm8bc74EJ2OFcfPOqfaF94nkzVJUNTx7XADOwac+sASPdoNB++SbLF1
/XWNjHA+UABaHWmjeoxfyMXmuOKCKYmPOzAr1HGE3ckX2huZMIdq0iG4vODoOQY6xFCCl/dQc0et
Tot2cMaHtdskJWZ+gEwXHindvM6zEZfuhBiIH0O4eg+jTBCWw/V/grumdVSRRM2/m3mTgJ3DRWOB
Ko3gPQztPCr4pvZh3MfwQRYmJrTji32XbDrntAe+P6u88rQjqPQaX58+QsT2C5zLTpWlTEDqBdoM
zjXuzIrTQ5p1gw1QCwKnfBnA3bY3OuErQ59x/3awOR5cPHVaq6+8liveq/g+NCdLc2nVRiDPyKOJ
dJscCotV8lwMJ5pSZZLlGxFQrMzhxNRYOUDSUIPOuYBO17HLVkZxqijLNOEHurd8RVrkHt3YAMDU
BAWgunsviUBZq1Xwu7JCJ5V3OxOYsBIE8rwPMDDILUMBe009RQtq/otkSEJx6iIdD2QJF+ieXuPC
19wZM/kB9sQwG1uPlE9z8yjFBviZAXAl4WzZSKtVouI3cRKp2uRifn371EXxKvQD3HpcPSbPVLfu
+63jZP/CPLLtg9CQumKmYOBgFU8k6gz5SVUKSKFpny8NoOZVlOccImbvOFCJzvZ3bTUII2qmvDZl
lGrC8zqdhol87YXcQWk09BdUq0P/9O+IHGGh8bsqMSY5632/CE4STrUy+0ICAhKdeUDNjN+blXWZ
Xeju7w1ZAt00FbAqoRzwKInv0YgNzG1q8WvTAUN1D8CFmDDtSG2A056iaxIzmfJne2K0+NkroTi8
o7szkO5oIevWX/++dYIEzAXwfWVznsowQYZpLrslPL6Skc63oj/pMOa5ctYpprWeniwGnnX59hCu
PUHyHmKUGcuSiNdAD5hrBeXEkBWi3hwoesyBn9a2UTBFN+bBRStdHMp0a+nUvIw6e0Trzxby7ret
cJEpp7doMNshe4uWUDpiwzFA6b0TQoj725aJi4xHiTEeZTysyiIRHkKAkk0T8oeCLqF6NJf9F2/M
63cC8OE8D2OqlP8/ixSSxRD1buQcuKaOjLK84SlD1/k1tUtQlQ6WYOBUN3pcmk76EvwcLD/g7Uzp
L3Y/7komyrXIPlhbNK/E+5IlaV13DWqB/A/EHWYF83H9/Hdnbi7doMfcKFwHgIYzyVpIjxdHx15I
FYGzhFkMShQkpQOUvE6eWwkizC+kxrkdN3p+5T0ZlgSI+REZrS3aBUdEDcMuLPpqcOzmuwlrlh7a
NiARLmB8nAbTyeSAp3rJIBL5ejjaXw2y6RVl6JGfKe2PIMNvmMbACzGvu04005T8FiP/W64C3uAe
Fz8yMYwMmXtSYm3uQgFofDhaB/mM0y+lghX6B5fli3qJE0QdVeRu3g+fGJCKJCKF7VLdgr7oE1pZ
20qZwL73Z8qopurzrCUI2jyM4EBIWx/FW2Ei+ElkH9zMxUjIMR48lurIFNQtk1kkEl3T8VSwktS8
VmigFw5HhyHH2uxqEGxXTVXrChsHUHWSrM7i+eYSqJcalFLD+uIaLtkvSIvo6uS0AsQY5qUwRRFm
UOTGlWQYlrT+eMi8pMDETjJWyPdz2DUHMauHe5RrXhR2K1LYtKO1M95sFbkjd4NZw9xYi7xl1enZ
DHM8l656Ey+CA3pz13ZEfMgxc1LRsAoaTaLqS2ybxsv4uEhSHrWvouoaso41s4RrFqaXaK1/PqP8
EefJMulquau+UBEPDYXS7KOr601aQiM+CAeQMYs5vew9sTfLkIthje0CJB+VkXVBaF+yJt6tazvF
cE/IrT8XuFILoe+27la+M0yRzo3/dcmbCkIjyaUTu5TFI9UPshqJqCSNg+ryvCQW9+odHq003onn
LrI2JPWYXFkJJ1xTVg5m5mbQIXx+aTIJrOAoWpgdCu8UbUylSYNfXLbiJDh1TPSuAWPad4qF9Ri4
VZuiZFQ+J64k2olpsiG6BtAGLV5M0S/z/IBigGdOHyahZ3kEvJaI2cMFRNfauivhZPFUqktk8Nl+
YZdfse3ZVIt6X7HhNXWZ7mYJ+A0efCf3ovF5CqAIwDtKJ3skEc9dLd+w/X8YoKcV2hfm2T5zZD5Y
jZt41w1QLEwcTxRnKZI/1qwMk1WWiY0U+g0B5EmXOC8oV/QaxeU8+0kqdPqL2ZQjzIrEIloti1kt
IHDCYespIrRiFf9BiTn0RKzHZLsjDIngfWS2wC0kk6vRnnphGIiKDAlmmOXrNTys1FVZfyENCbAT
8NEN4pAJ/nrUUzffujy0N/YRH44be98skPuh4UT29gVkyG7NUuo+pPOhjm8Gr4JvIfB3oDyRlr2V
xwfNaCcSwfrXPcyPrDaHt5qgHTGdrlHbqx+b95my+KjvLjSyc3InuLnGc1OgXUbDUDAayHt9SfUn
7uoq7pVO+hcIM0WwYUNLkCC8GvicM6vag6vNSbubSgaOWqpJOJB2J1myMK+2THGJH+PLOxz50woH
IqegvP2S3N83MBMMgwPrbFrpbixCQQEniYp+uIuFJPPy9Ra/hpXStNI5McZw+A9hCTVNcfC8UMDN
Ljj/XSEXZOGv/Ttqe1E4LmhKqzZB/MBCvST2uM2doLoOra5N8J1XFNd/NWm+WnfCtICRJ8hl4Emg
81t08Bcw+Of/OLLFG2LR0vkgi3p9M2jZmTMwwKZeQ+on/j8HAkd9Vnueaf3OP9IDEr2oU8Ac1MIa
dKXgcsKXcuGsMT1jS+/ZWix5IAby24VWHAEStuZ/LcMIcxOjn3SqXMHyp264R05e4mZ0xnxBBDvd
mZLbbynAihxe4taUATStZNiUnlL3J2QaF6DeNc/FbVdIkAw8ggh10dhKpKvcAFaTNRew1Fz9rB79
pVE43OYfyB3dvZo4URWR6xQiArz0QnFGFHolDccPTiJsQyz1unDXQcPK79qAHUN0ttVXGA0Q4Tki
wciiy2kmgraJHbuuaKT1vHshLMVha7u/Nm4NbqJ2hzFvicmNBPu0rv6CIDgq7puplSAdp4ApEuEK
3PUTCagiWT50JwacEJurq+bLUeYSm6j58ulgnTRVWc9M94SbXt5Fqpdx91H8ljumraF9PThx9zKb
A4Xfba3HSdDmsAt6N1Vp8r4wNu0DwNYWIUUKay2IQLfOTMycBez3UiRgGjfTNOUVb7tVP45CwXsy
O0hDYnQXF/uJr6kk+W6GpMMvlULwaNIP0JS+TbAVVhmhoov0V0Ed9C13lt0VuWaRmo0MjY8Q8f7K
KDJRUFwRLe8KRtFf+FGHMAUi9zyYvNKcpfncQeFTuNl7MP+NUnAHnDrApcyKJAeHHvlkB4zqlebX
/gL8PFhJm12X0UVQnKiVGSku9VHZd+5YXFojRVMUWXHhAYTzfXtZcwnP3wvCw+Lrwl779qbVgUfs
XdN8bUb8Q23//GDEKE6n+r7IkVDmTKY5rFi9oXC700bjGYLNDpsp9UwNaDevZt3rJ3cWP7HSTy49
C7ZyD4sk4fnlzZpAVPBgXUMaiPb3XYqMx4KmaOjLwd3CUM3h0MIaUa03ffRx1t6lr2KgT5OAjEkS
DxcxWiWnnniRG7d+tOIDvkJDIXEJKSzU6SdcSj8aI6Co8mzlhLtZh7MG85U7ady1a2+L0EtQYzGj
ox6iLRBQxW8vlLji/LK1BX6pcH6iX35nNmnJ1EaIw4GFAdVnv9kOQkJCO4Y0zZ7QYO0hox3vDzLL
aoZVgGp6Qkp9YLpRhb1tLhZk21nt3yZOrORGV3I5Mf19Gt7ufU3UYPWsx3ajyhho4miGtkhFqXuS
Jp1EhUi7FveN9J0NriubfAq3tUD2r05AEKCjttF9mTZd9iWL21DPRVJ3xMdo4VjAz4WbJa5m1bL2
U1TQFYIvLq0C52VFvLQQ3rXSFhgYTn7SQExuKU8sjZVrO7MF37KPFJ141+cuf1FnBYueZEffFpe2
ivRL6A0cRt6dkJ+YcOQqTc79RacjSNJAA18B6zfHJRG3BRJDTWx/e+X6D2hlA63Ho/cPSj5Gdn4r
PuezXXIxJ+Q5c8kuGTlmkIbat4s4zmUgkoaGsdcGxsovH+dHo9Fr5gZ+5Le3OkwYE69QaW0JqNWZ
n4uGHNXBwgXIbThv0JoRFDwiQTk97B2Usd5ELUpRS2IDu7zlCpKxS/+hxin6Cg/qQW8UmawqSOBT
Jg0HxvGYY0B2w0V7i3xJuy/MgbPwkjdtDqxzusQbzlbH/XjKC449nmc8E7DbbtchzpTfFnIwmuXm
VK/wIgLifJ5pJWhcveWgH4mxhMBnaIPgKCEp8PKhi4Dl7pQFZHohZg6MmeO8FwipX6Y0Aog/s6fr
2SsqWbazyBdJkKUPP3aGjGLxBiiC5QmTB+sIgveLonWGCvaXlUR53XPb24DbK/2ucf8rQDzVRMMl
/DTi76WWTw7mzYOqFGrgtHaFUdqqcyRYOx01nmZBhT8q6WrZw68mW9eb4i15W6NPrIAhEs5Eb8qr
tLvgxxktSSFv+kvvXYAh1L5D2Igz95cheeXeGisTWVtD6v7MlUtrOPp4SyJswJeL+0+z+T8gqWf+
BT9gPd496IBf3pVJkSpUjZtxsSFzKk0y+5Gs6g77tFNROPaxEswYnV9wJgsW+US+p7CMX2KvyJY3
vaCKPKOrGfEswkPOK9YKpIS7J54y3zHrwKlko8EkGGqp+QuCPryuiwpabdcIMyaVtffzbXOxWZy7
sYuslLzNJ5ZOkRCmP2rcqEF6MpS05TuPrS5uXuT1mC5VJNxC8Qghydl/wbAQju8RAORnv+MDXvIE
rLSAq5eeZRzLP/zkwkUH3frl+TyljjF3BQACoFWLDcnCjnzqqszYuoAuLiWkdRIOsvBzb6UIO4j6
MkeQHwLX9TWZD70WYsBu4cebWPtLs0He6Xt4s0PygjgcCOklf2sMbu0OY4xVTNxSugZfdCNbCKU7
mAV4IMnnjuQ0a8bvKqNuNmAxfLS3R6rwMRadrYOPnnnkqj12GyTJ98Rbi28iL4Ixv1qikGWSy4GN
PQ/8kgBBjXuFbIoclWns+SL3nOf72ax4vlAKx+KhDWYdC+99ARYVkKpaOGZh2y/tsYL9bYPms0C1
cDOOhQsV2n8D0Q1Cre+suSMdr5aEg+zPBrzQ/JlxUsQdxQLGQRQC98U9k9lQfYQv5VU0oRJZSYCT
vQBvehMCE6Hj0H7lpZYVVSmyVUxza55Xxddc/218G0hWkdJemvGvZdMtFZs1lgFWG6SGnW0YN4wk
+df6EnZle6CQbQ8v+gjOVpKqRw6HdxtT/+cAD3bHNFxkbM9zkeSbCkRp1Q0PD/5lTJ4nnoVJVBDV
np63m83KISknQFMp3hSM+koAZCkGvSh8wWQi1YLNuyPzfPcAdVPUNPG6fKTmh2gLa00ealIkQpiK
+z/uMlFVZBbEeLHIhT+fG/YBQWINEquT7MVJ+tCstHC8DfaOXLFSCdDx/HSOvCMVMDZryY6r5b53
VwhFsDCryPyPYVd8JP0LQz1d4GpZdY9GMFQMLtAd3LOxsPfdMjzSgZrDGRE0gJYT0gu9mZh9Btm+
2lp6RiKnV2Csag9IXtZO818fLQghqgkK1AazOZrEksyPw+eDF752zZF085o/wxsZsfMfoMHEhnkh
XV5/ICZKu8CnqBoszrjwsIfVn9sax6K3lh3UmQ0PWc7lQGOyw1Nlim6JuDHj31kSOguBDNJwxarl
BVcCU21xZMLttP8rphzYzT1EDDreyYmtVGXGTqgZAR67kI1R5DCozFhZvrO/8liNVlhwMZca1Ne2
EWiSWPYI+3fRPXBANuy9+Vb8NCUY+BAwVSnHk2qCdcGOxOc2CPIzoa2vlZdyCE3RWmnB73oWVunT
QzRbbnUAzzWZPX6uWldJ45VOn52F1KZ4mDszD8deo/yddSB4d/wAjvhxJoQfo9/SoCxiJbE6hYOH
Vulyzayd4HgCzekYC80Mr+mDSFyajDzIJjZtJ8GvIqtpNdvMHO4CInyXSgeHylTX68aqJkjwrXOF
be318PEDx8H1c7/8ZXdzp5oDN22R7xeDRWPGg4J+IHM4CNgUWRklEuor0cm4JH7ZJXQ1GM01ieKv
vK60fBJ4vI+NZer3gvjfZFtsUMHB+Ptmj9P2IrUgYQD+5gro95r6iPx8fGW5bXyjquZuRgMellS8
etDFat7HCN+G7Klam33lg0xp4uIgRz1SCDDvtljRO3YF7Xv0wevf5NImV2vmg46aoy2FVuP6DJzJ
0xiNoiiAln5HfkCmA+vIsAZSj54Fr8hYUI3y3dwWMprQHsMsKB+zsCazZxEZJxZ5bcYNBIYLuoEI
tEl3/zH8f7AW61JzvwTxlvPdnV1LAKuQy+VZQ5gQRulOtScGHR28NiG5jSRWZDGjqzw4/jMqThDZ
r+cFOA45/s52/E4NiO7ubL7edtIYxa06dTyh7XqCeg6y5urdRAgpGU3MXfFH/Tdwr+Y5YndeoRCs
Vza3nhYxHPanS2CqcQE9fVwpXFXZIqH1JePVISwv0Xp8c2/AqO+3HUy7KQyCHN5wd7NLt/X4NB9c
z0LveRmIBMKQZUXErY45TL82cUNDDFMoUpGvoNBpcVw3pnsyF8+AbylywOaYKXl+xgY1CflhQR8N
Paq3Z7koYuaCFowEwKvtLXk/pdTixbEU3B1StPLKum/SMEGqwnCiwRTOvmrxVQZwV07p6LFX/YlB
wnjI2Ey0bVXCwDQz5Y3flmaeKRCG2YMRZKDk2qXkZGuEBcAelbiqrlHlS5j4sE062p+aR1+rOBu6
+6Kgs4Y63u7+OOssnMbDQDGU/4zt19wDzok+oRNpyEGDPeMnbkz4V6gsLv5IqFb2tBqL8ZUQJGkM
8nWY1WeDn8xae6OXxq+osJ8NBXpVHfB5aMEoX/DDbrTdcMiyuAd1cX5QZMaa/25KCKdmRrK4MpLb
yY81J4Qol1y5CClgTRPcI0Sxub4jVIcQTffRlcN54AG2v+qFavxQ2V7l80oaH0XBRMM+0/HwUZyO
phG0RwbajDuimpY8H3hwnN7UBe3IXL/xlBYQoMpe8gtC8e0Lj01evy5oxVpJj3/evel2sReZkl7k
sxv2G8iXFZBbzMnUbKJH0vc4tmRLx1v9egneA1rUyaYz/vxccZqr0AtfZlnimj4+BoluBjdpSk/V
rM6SGw6s7aRQtgzyKHFAwZkDqIo34aki7fBtOPCJm8dixq4HRiRSqBMQR0GLEHfDSb9iMkhJNtAs
lItIkNWR0iPeRZO6Nlx0iLcFLSw0LqE6iQxne0yDbhrmwfOxtHk6842ki8X3DhbDeKZ9iUzAWnnH
hF+EQLVFqteMUBfWFJpauOWS2fPhnyvcFUz3hjqfaT/57+3oKNYUMkBxlZVj/hhnrooN6XQIZnQT
0ilvgOhI7OPsSjb2f6mzfelGndHOtlXaNb0zh3YJA70JGaPeJMxqFVKTKgxSHsvq4RZD8dLI0cAV
VVXZIxZvk4cc2oiP0ETF8DMxF7zHXLGB4aBUm+MZMPpYq24agOQZHMX9iC2nF/nFouCZHsr1XJxk
qzEWdOR4viMuBo+eKg3EzDZtXT04CWoYMyXAvZurBAuuDySZcM/t+AR9msFTmjTu6F8ofp7pCIwe
ot5mFJbzys7mjAGMrlTFO5r6HKq7eAdCN9D1ewvlPve814G8qMMMNbHgc9RK6jy8NKLaZlI9Lw2A
wIzekrhM4363ep9UgyghJtpfnep+eMev/CK5pYJGtneyRAEjL7XWW3u42qpDJOcwibGDeTLplqwP
DEmAHH2phUF0DiXhYywJUyjl3JOK2AECzHnPNJUvk8/wXp5u7zvqL6kCaav9sNIoWYIbECGhFkSs
N5l2kSYTiadGj5mPFqA2VH0qj9pZVwgH+knsJSjFO3EP601gNCDiTQPDgmVoOcmkAOGYRUlGgH8o
jVGc8IvFKUIWqC3NJHJok8vawB9Yf3ZXtcIdyBvz7H0YtvhIntSeTyzOaLybZp/NcHD2qMqzitmU
IK+XtBX9ceFv73ucfrR341TPIBCV+Kgl9YmCLCaCDFKsX1HHztPS5h0Sjpvcq4DUf8WQOpu7Q0YW
zlm/uq3UMsbpjJXmhS6dbDswLD3yZVYdfKRdbiT5yBvQGbOBGVPudN/wsmZ03B8eW86KlfNnRCTZ
6uC4srsIlLp+wIUsxVuDibHnMpD48bmF9myaWj7W/8gBUiiFFlUyfjIM43wtpfx1GbK8pQU2MXMt
BXXxprqREdcNlrH9ShZaygaUlfyxs8M6uFkQBidzQvUz6PkOcGVr6vczgp/qHzv35FhGAOKA1jnA
wOoCAgxKNQWJWjxoujuv9RgYTEik6k+d1Ro1KRgkAEHBs7RrH0NoPY1opMu6xaWk4zfS5GCl3PCc
iYgWkSKk9gdP2B+2g84g1D63rodbBzthYm2gCO1Wo8aJzXtmtaJFfTg8IHs8a8hAQHVv1q0FZfU7
vCidusgsHlw6xfM8IInLe0HhQ/1QGaRD9MpfX+ouRonqlUExTVthT6fwGXSxikb94pBML+5Rb0wl
sk6m9/gmpSllQGaaDyyP7peqv51v5nIKjk8mjiUV0jiLOsEvqEyQajrpIFv7Guhi6aKbK+VeZc/6
/CQkSDr69Wa5oytMFtHgAKz4GqNXzGEA2oRcfncgN7M92rq+D37ecs7n0LUooSnEQJujpsd0+NcI
vfGTM5VjRMb69JULiDURSuF0Gb9eRiey0vbcebfEm0QdZt4bI6CcgLfiRJXhtVlLyGBvjzbRAeI5
t00MG1JGzI4OPqhJdTnenAzfGLMofDscTwOy/VaWbMJsC4WQJwO0Qs0XQlg8j+wDtXR12Z8jyd8/
vQmMeBuXeo1T/ClwQwKoVNByJLtkbUbhE5C4mHOPSx7e4LTA/EiiQuuBEThoMAlYRx8cAgZvnbeM
VJ7+rJB0MQmlfNWNlDjkuk2jVuUtTCUtHpfphNnzbclKNyOulh1XNFspRtssuq98b4qiXT1W5MUo
cM3zRQL47xC1k7svnRlWbuQdydOp/8aVXVUDBlkiy5dqw7G0P35kUc+uvwYlIqP8AQwA2p3u+B3p
qk+wpiDRK9OISN61EktWrBgao+ALyVXS+Kd5xzfpX2BvTJjJqimWtczgLJpz1A639s7J6nyVZGdF
eXIa/sMrgjfj0SoJB7xDYGZPwgv4Aaq2zIyhUDt1RpdUMgfbHcrUhuRRqnUDq4I7HaRS3aph3VwW
ttr8ybHWT9a2/OJPL4xXfsK20tZuxOOGrXnaF6II1p+bJ86FXs9rai+kHMKmrqvrIUuQ3x/oDRH4
WIO6h3KHVj4VV4CkcPGYhroYLLxHBmBQN/uHIiLyElQZ+NXQWAlcUtru1xcTGQhDu3mQTIbv8J/L
4hZge56i4F1L9sTKuVjvc1sfR3sP2N6azEXyfD8fAf9rSQAmNWzfq1Sg68IuJHV5xn4L9qPr1TA1
+XBwfCg/OzdRudUYFh3cjce+x2WT/CedSlmx5BUUCEKM4hqko285YQJI6ab9ZQdAx0RRIjiafO6Z
LW7354ecnQldzqmFYZdjYHOIc5OX5pKs0NX0Is1IIj0d2KOPxMCZJStVIWrrZPwoRGJOSINHhPO4
SxZjkaZbuXodoMUviBv3xqDaG/BY5sfENxe18bdxViAEoehcKWHJ8Ra5aaIuC8A54dWD/IdGq0/X
PZudg60DdVuGUh2BT+GYDRwSZKpBpYyYPifAldAKEp+X4b+mtBHoUSIhIiT9eKpTyvRQlyNkCFTR
NgMasC2etiGKr3VtOSa5mcJoTRnsH2gl61RLe04c2z4L7PNEpRDZXi2yTLJ6m5x08nF+HR0i6/qW
u4ugutOi2QEMSOJbcAY3DlInUeo8og0rw6qKg4OZ82lfIO/WnECVVAhZryGtCpm6w+asdKHxIis9
1neloWwvapj0dHnPk30HxALiLAhXn9doYsaYarIAa9+5wWSOa73eTdkmPgydHZ21Er1eh205RKp8
gEma
`pragma protect end_protected
