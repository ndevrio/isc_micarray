// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
L5jUu2oAX4hzUF4eMfzHdx39MvvM0uCbDjnLQLNWLtpftnznrE7A3JBo9sM7YUpq
Z3jSmT4hjUdLYN0vGiWaAzy7T+cThMMRL6u4XimZkbNkv7fBh63Ba+83yncEzgzH
FsP3JKTNBHhrE7DDOps2lyyrEHePz2YlAhCct38XszZOh59AoJXZrw==
//pragma protect end_key_block
//pragma protect digest_block
hYYjpKCsGrqtLOFFhJOoKZe+aH8=
//pragma protect end_digest_block
//pragma protect data_block
FUemBimcyihF7nFotxjx4vdv7E2TS+Wr1zO5RNVrQFhSi/jE+L1feXM0I5ZIUGEq
ds7LpiFFSyCMUCu6m9VJk+TvB1t2J6z2MMmE4EjKwMMTM4lZ0/dkMeLAc9hyc04L
58KI+F4VT2IpFqtKQBLWHoHHCckupgLP/0lxO1H6eK3AaemLfQ3oN5A+zKyh9PAh
dXqHu825cUGKFxiKDoxm56GqlDFniElbEMej7dL4At/5oesKUu2bjesU33IVsUhB
zKw71Nt7sQlKBzGPzeeakjmTM+7l4lzMezAqpPKXm5Cuty+U1B+3jsggX1eTO8cY
/o7M6+rZwisFuyQvsyC7PGayd15mLhV8Ec0Asebe6pFwBZNoN5gwywr+BBpYzPoL
vpqept7IFd+nrlGybsVxu1E+NSL2JoKD5ipAGCMvr0cb59ci7U0nLq7fMvQR5dxG
fS0nNigaQlYoKA3JxgPADniLzw3Lwt8DqkJm/WGwyVDzpr6891IfbAg1Ub3r6D7g
2NKHAWCTl4lbpEBW3AAMrFUpY0uB5+EuvHm/wiCP00Y/QqKWpvgqyxpqq52kSNCl
DKR9aSBSYwHIgNgT8roXx1aG1VCJWs+hYaflQkwQOdyOuuAvXi2TfQ53ym7KYldT
7mj5fMzsM43Oouw5L0q73QDNCoLjEp4MLn8m2hHLq1KMB610GcnWzwnTaYh6OGQ8
hELZoihRkydc9ryuh7xBwYzj2gFDQltF5RmfWpfcQ0lVSU8ZJg4d6ww4NdtE7JJE
buadYi9hXgQvlc4fGwE83mxVBCMxmlYfCdSPbQg+NHIGh5LrqPOfIVDpG/P9Y9dJ
0ic3oNbHB6CZAVSVKEbad4Ff+FJVqK4XSe9dLP0c5+suGbxZJEzg3ZxxaI8xePza
0f4OKVE6vwHcOQf0qMlZY1puMv5NS7CVcymp1ATon0NHnI81AsTlY2DQRGP4RdwB
+aEd9ArvpISIPp5ToUsBaMQcRFNWVbnVzXzmIhcijDXsVJO0u8rJg2wpCCKt0mW2
phmQmBmBoqz/zLJaX/wwcrTY30CIGm4GKEuVWSaiGk5rX/n6DOeRbKmAyczrXClY
oicDumIiEYG02+XdAA2+B15ucMBOxjSwT4HGBfNRJGn6pLyz2LasmIFABwrYEzQQ
cj52ZZg66RDXZJ39siZju9CmNmmfiIjeYrWu/3oLO//XN53fNXAk0+fM5AA/h90/
Smt2juU1KQ9+jIZsWUfiFHTxQFdNmRc4sWlUJDqsdjwHx8XA1QBFJ+msnozB7C93
Kbs6JDiEjEv/7iftH05OsZtBmXTxTfLUuXc7rhGn36pGIlY6OehL/MZ6PKhEd7AH
m1D9F1oPTkRGGSFQNyhvRW85cHJo5dQSTHG8teeVBAZRyFrZ7vDGc42I9IKF+9qc
TfzjWj6hl1P5KJtsHk1kbky3BVAY3HPEubHKwUj8A0J5EJLC5d3EPDDiU9RG6i0B
8YWWxl0Jbrbq0exoXkV7vwSvgaU9Bkvng89aNv6Vb0FglzQhB96ROnGw0U1I7Cbh
G3JuG4wjzS70r5+uW7gE8Sj4cMcTCahxNjmCfV8/M05z4DJZ8cv3qjhF5ZV5aygd
tkFs2cyyNP3mLnt5keCW5/dNOK+7UEA1r3n5bwKQZAkVu2+BxXAATRgE26fagn6r
WkJYydJWY9CI5iVvsKcCE0HDpWHYvd/A47lH1+72gQF8vIlevIFkEdarqB4aoBhn
R16AcKqPSBuiOzqQg0nnY4S35uXbG2NN9k/EHtwyaiD3ergP9Z4LTgI9JwoTuN/L
H6fcqiXF0SCKV6yPHOJI99g3mtcS55KqJo5LnptPMOMRLTrABrcs1u/LDdyZ6jQt
iB/FYa2jyFCEU1sTakCV074hbhTAHQV8ZfnWFb434A1TknZLfU9mS9+uqidS25qY
WihvYEpxAf6+aBw2NnQNR5In7FWBqY+WIWpJ2jcB5DiR2fi6VvyZ5Ep+daJUlHMp
YDULn0Dg+K6fT1gdJdU4rqDKzt3MaAn1oqopTMmjLzWAyJTH4aQiWRuAzngirc5C
mwzL9Xf97kN6wlPf0vh0pekskByFi+00zbh/AKkl26WiiUTKAjos6Af+R3uYw6ON
SD/jLNl9RjxauSDYHHPAtMDp+p9eoqeJfN3fe7a35DrSfaWA6ixv3O7gdhPZn0SI
y7hC3Hw9lWPYEIYoj/Nk/FSCsf46ajnNuzSfSsZts80OLg4C30ETSnJoUYTaRuQI
+5TFhynqvoZoCOkCNuSVW3Bn/d1h8U32GLsnvJUc+WLk3AjGII4yrp97idTJhQXU
Ie2cqFxAnBc7OLClnUxjazkaaNaad75yjcIYbfamXJP3GsNgKOwjkAYC16U+Y9eL
EzXyya9NCLntcLwotcHlfjVjiHimLGKUe0gCR6Fg1q6CWjck6OYnT4liZdsFe1Ap
OzUqloULWdN4cJTmQODN1MxPfZWW7FtLOlYfQcNopOmebXepw5rbH+Z/4ivZ18vm
RIg8xRdhrgP+dHu+4cjpHOZMj/e0OR3I9rIbSP4QidSQppU3qy3O1cVeovJN03Wo
oeJHiaPbJ2cSCJMV6+4fdvuwHuiWJlC0bNopnuRV3e5QpDDEb/j0fqb5uh4KZ/YP
XqqG1KIf+tikwdFyQXBKBtDeilZ5V39GFMtPA4nRqIa1OqgihDN08CQCqtSOdrEI
zPPxrKcmDScB2Jb7nP5TJnzGP1ElNN/6FQlEcTnHQJIXTLqfkH7nkNR0ppsaWb6B
iTVCpVyW7pYrbiMK7LJAtAP85TrqhV9zv1mFF7BE7/OXdLgF38dHFJlPxAuQc9ZH
1r3Qk5E0pjVCk6vdL2XFoMnlBx6+KxeUwsqAYxeuTKNWrxc+R3wjpqAVgpkCNQup
1a67BUekQmY4asI66qQSfANWjeLK1lKyVSA5eM40sANlKYYRA16i2UzSR4hOMKqP
EGl5K55yX3T6gxvF8UrcLt93R5R1uxHK/rhkz7IiLeT/x3U6noCcizcnWSNX5D6q
IytlxyQjHd4Ta1RXUT5QBrNC7ANqRwq37ca32Sbx2iE2TwVx2MnoGfQZ9FRgOks+
WmQA1+Y25EZVZ3ZB57osZsv0CeAZaSORJqA99LMYmgg87GCZ57XfQOmiyiEfUtK4
UFNhEGFtxDXC246EAG6M3GAJiwwPwYoRf5LANB6xCECBSaUyV4GavDxzEw7Bt3tA
dW5XB27ah0g1AGVzO0/2r+dBCnZ1zuNxM1wgw+oJrbRjwWG9OKGpnXr4d12zu5uc
/gEJ0xsrN447FOPd5aCSQA7uiJEsbEg/6SRyfrR05Aoj9pGS0ROqLqkmr8fr2Fhg
LxupLdPPdySo5Z2RbxdG/pj1BHrqwYxrM9ZZ8RpZ8YDJGClQQpDKYljjUR/eL75k
xh0JE7FjzAJv7cdm3ECFe3CR1QwIyyrN1w3wVLDx3cGmW+AONb6ZbgicoTmDgzE9
aQTTNrbXovfMS/Yw7p+KJ+19a7DcWgr2Ex1kJ1rCy8B4w8HW8S7/oTNhQCYXOt6b
AwR5r6q3SDsz25JTbV6wqlJfYRQxhK0NoZ3LSx3Uqg5wNlFHiQ012ScfJlM4dWuj
zjLS4LLUneK294WnbGaDRRHApfY2PYuHSNWqomDvIHmmt/u63HmDG8UnrhM7QPPF
289TMWTWnfH7328TZAbCt7fkMC0P0ZDBtAfpHoFmh0R/DewekQXOsaSfm6KV+9B1
sMSo4Ukc16cvc1Xexy7vw6CyY85Vshdu+n4dbVxZLwQpK9m0wsmFVPJ9kBGAUPJl
6btvDg2vR7G6GeEaN+SL+kP1BwRmhCdeVGyni7ICVBQN7S4HlpxxsOunb4q5aV8Y
ZtikK2uj81JQmN92xJD1wOBfy1doq9ecq0qdT9H+IFkXO7ji8Zgju0OXzsg18t2q
uQp8lbWwzk/cFobICexT3jcjtwtYh3SR9a0Dr8eztBtbbD7yjxSABanXU4RaziQC
KmIs1FjRFTZ23tH50ZU1IfSh4hAp/fLQGJ5iFE+Fk/5OJzxNW7LNK30rPFGIGG91
jp4gZ3oJO3QhlyNbHjihpD3QcETXY8RXhdtWXgWwcx4Vc5CeiHxKy+tEJC0NvY36
oZHI8zQb/61QoqRo/M1H5bTuK9KzjihJt563rUnjGagiDtgdOolVQ4JnHuV/eQiO
dQACQ83+5zDj+Vl/b6AVaTPB79F23akFKAEEtEAdPbZe/Kz+WWCWL2lEGXG7kH3F
T22NuD1B877c1VU9Y19B/QRkJ6i63/Xc3RgXRlXtaP+qizHjLaYfgaGlO4HqZBFS
elpeBJOIzqbQwMe8meAKnbuzPYh10o578LNnQaVAsDQW0PQk2lAOBLYYR73zG+gI
nDObyT8zuz00k18+JN5ivizm4t7cY9/v7re/3Bzs+9QX6ReI5X8Tz2f74N2dW6El
CbbZsA+zofjTjTvHgyrBkI2aNFvz147d5j+gIM1Nwbmr491nhtVBK7ha/Y1moIz3
NJfHfLv/mP37g2cL+ITxnnMCi3meqbq0LwCUwgK1mwgHwjHNuJXYT7PQs+senmI+
cNi7R/QZFmPKZk2d88aRIBQlPbQt/PLWbmX6AAYKs/TZp0qClwIT7BKIN+oM8Mpw
phBE3XLre3MXolAcM8ctbkcTVnH/alOy6e7wnD4fbir7IeQRqQ928q2XTA3YJ6sq
cQc0FM/7oSFL0NMV/harrDadSZKLVXRMSTiGtlS2R3N82LTDN0vLqBT4HzLz/ARY
qTgus0M9XQ61qf9ouM2SgigfsKNO1xK11i+Bn7PNwVUFiiXWj/QLbBT/6DnA2JWg
hW1yPQYg4UnZ9cqLwqV4cZ/ggJMsoo2OoThkigt8IvkHpox+ktbmJByzhwPjJY6Y
rwjA6XFzkZ8IiFQnRi0hQHrnYxulhIvAaPOoAbYSs0d5Xiy4q3jC62drdUY7XPdc
f0euYMupeI/1OzlVK6nQV0DhhUl2jbUhoYEYPWLAYL8wV5KfWggQVNvBAUOnFlMF
OchZhepzAZho3Jw6rOcM0DH6iTqi1ejeZ9DGB2QFdZ6O0AOkpUaWqOseeqTS45X7
N1nkTzLiWg/4irGEW+77JUXvoby9zu2bR8qS9Z+Aw70hs2sDgTUZiBfPG/1HLNwi
+aqu7lM60Yi1yzb6qye7a8xW1+/FbPfU7XzoUa9NefQUsgKaWYuWjBqJS7DhHCbr
mqDrb0Nw4zX7DxbPeiC5qt5DdenlML2aDr4kB6XPS7qvXMvRY4NOAHKE7WHW64Jp
8XAdWZyFnpOpc/dppi/OGml10PvrLr+sIMMyTkFt0PYxGKZrXGFxKOdR9H3efyQ8
3xssLFAtprwauPOKOhsPmKMNdi/PBorO3c7+vUFlO8Hp94NwnbnDl/Fvtu2Lo/pi
wU8croIi1cbyPW3AnNeXrK2ptx+Tb3mNPQMbTJlZ0iB0jnbfz/IGCVpoR4iZAahf
cxb3sAI7laB9pT3CR2KBJoseisKkIrwi+Hz8FLZOEIQGl0qd0t/f859YrNZ6gTEq
GAVBRqFM6u4n8snayKWstlNkUpsXk3R1sQsjhfxyIDsN2mbEe8vQ8IxWCwQUrXk9
uIv1lQaZj6W7uZVIBJzAncf/IYWO8U9CGf3qEe0/uvFaM6fajuPndjRmbUc3jJGJ
Q3FbnKHaPXYN1I+oZZg9k9w4afZzngGJgWt2JftdpK+k/wPhs6JUDMX4YgFS5pWl
tRvvYtzoEATd6mpAX7ksJSp4b7o4T8N0r9K0A5H9pVeJX2ubfyxF4F1lUGWHxkyi
ELkyqgqZsCtz0peWt5BuCynbvHrxBAQaC3KTlpApEJKu5s8W3vreE9NtSBbwvkOr
8JnXjoUnlaWtcajN2W9mjTTmyEu8Ww+9tGEoS0kqkCziKtthIRcnF+IqH32Xrlya
CcJ98Xt0uOGpUXw9sEQVbHMDGf1FIT09F17ZmWbKpPNa19VXf8oVKbE3HmLKtSD8
+G+9BteEnbmAGLlEMjpjHd2Id2Y2hUlK3MMGCYRkL4PV2taYmjNmchyL1tLPDIU7
Jm+J0ZjD/9HsmzO6AJ+jHKIHct4d2QF9wwiklVVXAeHsaaQh7RRrbflO8dBX+TDm
mynp3A69TyECFJkG1qJL+rxhepGTJs3yb46JX5i0jOe5HRzFmvTscPnKoXUM8dAx
xncYhRT8wRnQwSTHKsD7DGgTYDWxMPhnjU0Y/OZmDBV3XENDEIMgUyyk5e7to2nn
CUqHMXeVpgR/gVNVN4Zqzsfq4cKrEcJdlSaJuoxl4GP81B36ivvComwgQcZIxGFe
ZTIw/eaQtz0uehZeHB8elnRvTfksDtLgh6K6Swb5/OyI7WSTSOzf35IKpx7Mrvlx
NwuhhRHHtXAsvBR0D5QlEYOSXP1ORtnbkzNfEwHfWJb4QagFTrmJ1dV3jorpuJy0
SW3rdSEjnWXScOqA3+1mDsUkS/BIgtVlCHo/VV4Iq3HQyclUF2+kcMPNnE2Kujwp
e3qqO8Fhw+UalBuVDmtPPg4sFdDl4b01Tn+PWJmyVAHZcTsZSBpLoHQYDPpNDK1W
LDUmXdb/Cj96i+7kx5nt/SKhl8QQp80zPaiyVeZ2+qOBf0IlqJWna6IQQdMOYQvb
CvxCCKNTC1Qx71yP4FD8SndWtQZ5N8n2triSVQLkr0f3t2UOzAiebSBMNM/b/GkD
wycyZJwy+4I3sbYFJ+/ql7QlH13jce7/yQfqcfdvE4/IOoyhJAh7KL+hX6y77JOn
5Cv0p2FUuM0imdAGyNMzwwo7Xys32dDoHL3XDyW3J+rPhntPVNZwbY8I26BGC6qD
n1crCGB76I4YEeUF7oLO3yrDoaXDiq17STA8RMmlGZCT2ksghton5HErTUIep0KV
QamXgk5CnCpgHLZoHFlnD4aLKlsngUBoU0S0StLEKHFXSasjxynVCM+icuO0hm1I
6phd5r6Sur3pRVOEPqk+ONXpjqUq7G7/13xaDabjLf7HLROzkfvQvgX97EOpX2UW
ozXy4BgqZttsSluXTbMgP65zBkseIy1izj1BG8T4qUWl8vWP6qAIpJHFI/XHb4KQ
a7EdJklkI6puxMPAnWf5ygf1kqqwyM9faig/ZsFNrR3H1I54qkXkWknlCEKUApHu
w0sV7eOg1fGxvHaEzofphsEXQGPSD5RgniVYsAypFzw24ugCq6U4kCSQc5SepssV
Bd+DWnlrqQJNgoYufjL8pLGjCPm9c7idQoZbh7U8VhM5+Z1ClVF1YaaNUiNRzoGC
aQJGg23417VCM6gdFRLFqLx6P3GneuxZp4+GtxR08hpWL9vQmnvpy420Op8GJFtK
SEVEw4uALpDNazy+J7xxSmvyxzSe83OusEkXEy548aB7o7BY+2HUBua05JGromI0
yuEoDueG+p+N56upstqHUjPgGaRdzMb/E3KkmO7Xj5jyTpK8hJrG2FkIbWfd6oCd
1nvkaf01mzbUzTOthnyp0R+8w43RGy0H4d41ibVnDm/SFFwt2mR8MfiYz597ziAG
Y/svmHODogBen/6QuXgbl9+rPvji5+iyUxEFrNiMVU84ALIlYCLcCfh3BmEhgZlt
DYUEuuxv7o1IaElaeX2Uh0fZBXluoDc58CoMa+9rAGIAJHkyyGDwLlOXzjDcK48C
wmQGP8CuvZm13MDJgEiINQKoYgMoyMHj3ybzn72lQuzWxvnUA3BtDc7jkpBduBCd
SvE7OVLU7qiiOgSAPz846z4M3VbWuKPiyLCWbxazrG2oVzLrQ5Ncq3TnKJ1JO61h
J9czsIhAT+U/h2LYwRrxapz+YzYK2nPJLCOuOe3PBXfGeEBhjzvkUIH2QW6V2EIH
Gv0M3VKZ51lqIiaSlYfcf1yoliT9ejYOXH3Xvyjk/0K2kE+5UGPr8N+i3umpysJt
MIsIZzBYBKt6uS44jHoe2aUNBguZyZZfKg+YFQB5uUpK7LZcXTmGvp9QnveNiUOe
5pyiBTqMM5f7SpYG5nII9hFnIdAhLY4tUTtumtk9QhTgHkYGYzwGk0yyVo9sTlHI
Ig8RO5rrIzQlpwm34vYkbgY/mTmNbquch+bRv/IO8Ylh2mGSPDocK4d7sc7iTr/U
3IQciyBZs9GmkhT8JhQA6kp/n+Sn8rEecy0HSdmnAvZT20nVoEIYVHr0s9DXoJCT
1Sk2C9v7PRC3zga6DXOjB9AL4/61gEtEzBtGGBee+PFfQwbCHY0qn3YXjHh8Gu/x
P4SanDFql3qzeG35zF8IinnM6yCNdE0ZyTg5qwHZFzSG44WezzFmJQl9tlQ1cjDy
E7XeWTJ+nNhCgTZ5NAPzRRVdvFIJPlCyPNenekDl49izg6RmwLylwQouHIxPeL7z
He9HPRKrXcLrn+hIGOlJI7cjlanSXvA9GYMKEiN0NGRgOoyPOggxtqm3pf6xvzAz
tHN2eBNWULeWmBVvWwppVEPtibtwUJsDCPJ1aben/aV4UO0OL38QzEyXo2S2bpew
Gjuzx7E/sjouh2SOZz8AI9FSlpr7bgdRMjnpJm+CanSxyHS475BF/z6bKwP1WO+3
7ZXxANKdoChNqi7p+W8UoCYwGKTVIXXcapwjBa/W+HmAHrkAQIeaU8UJhws783KM
mHGqI+/0CAZzV2lqETAoKWwFaFtpFuvcRX2toYggZvTAcH9BNJk3FqUMulN8hF+R
mX/0ib5bnEn75XLqAHuxRZCthr3s5KzGnUTLmhE3lZxkM+ih5s4W9Uf9fkpCoxp0
eXxQOY/k5r0OI1gWJgsuo0YQeb6HHtfofZn5Z6+u7/EcrvboApha9UasN4hpKiVs
Ampaq+dbe2BLkc5ZeRo6cJNjiatDJBaGH83x1aG9UOEBRGMN5PCEwChkTDqwR2nq
Z6s6xUy/6iVEmePGyzO9dJl357L9s1df2wq28aUKVaaIhPMvEaUy7mYsE2R3VTwi
1QZPs/4U2t+G+ZkyJvbQ7bxH2/sxKbFQTVuFX8KswfxYEx4h0wZtk79mS9fxJAYV
MLQdJBO5/6a+BJ2KeBzPprM7PDlkWs44UOmQy4K5Wtv2S72c8L3YndcCnXE+9ec4
ObQh9cIeolhto/637SgMTwIcV2EYiec2eDCkz2o1rjowsUT+cc6Kw+kC0el227HZ
Cv49siul0djyg1A+ERK6BturJFF+wdMVvuuO4TdPuZQDis1jOiRkbKT6TW2Xzvsg
tlb+53sIbIHW8ds3cO6nFx7prgzyAO0ifXz4TM8em4EY5W+8KfmODGEqeW94Q3X9
1TEPVACSERWqF86z5GGjNbjxccNxMsUl7hbAdwNEihkcIHfooisTPila0zNd0y6S
17XFdREPzn+xxTgSUsiP3JPh7Rseyfo+f8wqLMLjwexcQNHMKzI+LhqsfcX4tpoi
aekK7fJq2gK7lbOgt6iJl6Efh0LXKnK/tlElLeEioR38/Sm3g50bb/P2Mr50+fHe
cBwNWRAncXHmFFz6wLvDsvhBWA5L+77u4UFG/+BvLrXrn5fTsobXWOurkwI0vIf9
kqiPBKOrpjCHVQbWxTHHIKNzZESydiGp+khR2M/r/Yue0Q7bhzVBvtt6TBPZYbWC
9kK9lvWIjv7+tXUn2/AnUbKVg5IfRtRkDfdUpSuqOZ7444sNbo3ps1hNNpPSxLrl
AicN5arlqAD+Y6xP++sxXSIjAAK4xkPdAO27fx6K+zFA+4XvKQlwt8ptlLQRr6t1
cHEq308ywo7U+duWxyavv6nVIZCianoKIMQJhijOFuhHoiTBYIu6HDwRHmS4J4EX
eA4vwLMonOalVSoD4Yk+Mft2T5pKLmiq8QkAihHlKPwvEfbqIwfpe+xR3ZC2C3nO
Zhq6TSgrJ/vVNypYwXxYJ4aK6hQ6IOXBk2x3/AdUxfjQC+/bfzZsMq0waV1EPRBh
EpfZ3Zm62DjhZoVYBphbxnaCPaqEcxUyMCJzK0hlpONMyYzjnEo21iuoei6cqW66
hauX5hoPY1QfjH6CXM1iyMCDIUq4Zn/Ixia9YAXpChDu64bqv7acUF26T6ZtWB+U
SIreUStaW572D9mto3qkThMhzGcsY6dAV+pHEVrUln6UtQtqDbacGA+GmDzXvxLI
FCd5WPT7l9ZzMrQm9kXoUbJvUyrwanNsZg77hna7JWk/8iZ3p1HMaIzGF5cN99Mg
EZfuYakeB7zdAik+IZZK/jJR9K3jL+3NrgRlgJGv6pSRHV+hCVNinE/T/LRC9xw7
K5KGLUJL901pBqfTapWjEroHDT7Cf0Txa7G7fGdqfg/dhRZ0d95sa9/AvP9HDJyT
pSOkpgt0c59rZbgYHV749Ih1bSN7fHWJhcwWyFEPCaT6qyrp1FHW1vb+cf9uA/1Z
QOld6yq9BXsP1eBOOUloxRTb1nqonXE9YWQmlbMyZftu5oX7eOM9H87nrH0EKKzL
i2tew1uBqvyDn40xZEVz452+b7i/yYKdSyOscFVMpl6JD2yOQjFUdjLJSDkvPmyE
h+xwxbBYrHjucY3ZLC0FEBMQxysqSi/VZjZCdAhS8NoBuPGkl2QKm+cVZDaotuYd
zRv2Sn8bj4DhXQ0ADbEfPUFoORqV5OVmHj4HTONXs8NUEGfDP5UQ/pWGpjjnBwzq
6mZ6lDAhy0XG5T8mqFKXy2tSeozbV+ffV8/d52I49Qp+pRMuQ6lMWlF5UClySxDW
E5lHbNzPBKn0rxKfN6zKuJI3Mhb9ayJMIj1Uekuo3iJi31DLqaDfp9Ghv6gee1OM
BsYYSbSHW6ouZ5BdYFW30o+iCFaoOOlah/s29sqmwEET3yYCNnbjFul7YCbRGZvV
k6OsDpb9Ng1iEUp+nxfOEvwru+pcrhz7Kmq+isD/SHVocwFdO0DdSttvPqqWw++9
ytOxPQbTXx+P5fgIShm0UyRsC5pt2zA1IrTwRc9gdUJFgrJVDNg0oNRtuPfHlQV1
ycVkPKa0WLgfWMfqHa6XaR8sOW+daj/IjQUVwbEx5sRXPBZE+otjMSSEghgMj1mv
Cr1S3JcxBFr+XAOouivwcP39Oca78sRAZURdZ2EBVmj2u4qPMLM6gkxHYf84X6FG
Z4Hi4GGaDfWwe43BsFBdMBpEZImo0r0JTcNDsXTrqDG/dbtZR5PD39tORkQStaZ+
AUHpS/UuoV1CgK3zfe2FUhYj5tfCSCYLbSduPSDZnFlRsCLMFSxkXzZPWj7J3DZH
xxnRAPyGKjQgguszBa6AdKn4oDLegObHstB+eDT47nd3Vb3Ekr0ew2FDsyU1xJB+
zc8LbIxJUVpmmjI7kH4HITY+wEZAXM/W3nHYFl1+VAGoXhhP9Ys/b3ET9xD13yQn
7b6EMNSBm/c3akLOBjD+9OteB46iwrq/BBdZsFdxNBt5qiipol6ffaTGcHwP0sPz
k9lhiYOLFdqzWsD5z7L3GotN/3BEZkx/MiSSZbbWDjBUoxIxnhvc6/vXhbmyUTIV
uRmDSEDQ0Iod4Aw1WcZNe1Kv6Rm7lYzNIG/NwoTfF/cYYM3yhatbL7I5yvQ8Y0ij
/P/rWWi8LkJHwtYuuWiqf/ILuzHTmjAT9HNjFgv8Qopwrf41qw813E48EcUCoOQc
XLO6CZyBtuHuMQ7/TtK+1uPymCXZVgJSWfDkhdqV/DK1OWh5FUnsI78bvh2JBDM9
DpOjAx+KOYeblJuTCEdA+NqMvvLRrRUVl7cniYmSTdEN/6bQ+3Q3CWoTT/+Vp8y2
9sqx6hgljLng4unMUNl5sgoUsyw3P7bpj21iWKFI4yPraPjyoujkx2OTh5O0xJ4h
xftVHc9X8xs1b9ws+r2X5Pce/Llhe3sgrcPn63Fc3Q/R7CxeO4KQM/gF4HEM5mS1
iTEe11wjmEUFxiX2rzs78zDV6pyysJNe2Jx3E+qsTYXUzHocbyxPYYKCmz3IDxSn
UmeSgRzK2ti+wmJ4XX8B4Gkz+HTNGYZaj1C21lK75EUqQravjf0mW3BL3oAH7SaF
PNJDBqCERHv+/U6bo4nJpQRvPCqVKXVN0sOUqqn1cdRsOmVtM5Uy9AVGwnp4MMAt
Ws9IQ5WsXc07tP8UoY1G/MZQv4dPjEG06bpLEI9VlgBTueqj5q1QMuMBlMZlA9vC

//pragma protect end_data_block
//pragma protect digest_block
XGuiGDpqgkK/KzfS6c/8r2MGZ0E=
//pragma protect end_digest_block
//pragma protect end_protected
