-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
knxBqnGS7+9mdsJmjatFM094ZLZk8gXsdQI2cEC26YVXJaRxJXCdhSJ0fpH9SSEj
BzoGufR0LVo5GG/yfWiKWVnhB/+G6IgyHB0WAHj4TkR/D4RuiG6lULDtWlcRqFcF
P6eiYr+o8t5lFqhHBiqh4gsm6elNcreDX4Yl/BwkdzE=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5171)

`protect DATA_BLOCK
K9c5CluBp7eJOtqxBwMEIanImOACOek8RRlLjvRaujjw6OhHjNpQeLLWAzv25kAy
xJTTB757ai2AiBAtzIfKQln6mqAymmzjrNOfof/ZK/tmowXbU7/wh276msTR0VeC
Lteoi9ElBz8wBrTfAaivhbDeOSR1/fwIt5P0BXU7RNVaES4ZWuFIVCanP4EAPW4Z
e40bkim3/0EFRAwBB7qzLGAja15l3NwJcaPXt/MKg2scNEcNfuPlDXJ/5Xo6LmtL
WTgL4jb58B8yqf9i24ezl4InR8biXKnmIY43KtG5Ya+yZnotmlStBZAwQusYXyl3
9VfarqWoSS23dtqA+ZBRsJt7CBg0h0GZFwmfeCeC91IgM5EqPJITYK0UJYs0uvNT
i2+AxjwudieRFAbYHn5N+96CmXI2OrL6fgoKoZ4eNankyUpJbuyAyML6rG8r5ESu
22rnyH/hDmZDE609vj9+YxLa0c82FAPIH9QnzaFLTGG1itVBBExoObbfJ+jjpWuS
mzZaAAwlOcULrE+yBVT45D4Ff5HNhpEz37yNE7nHFKVGRV9/SAgFS97dTPSJD/1g
RuemmGiM3/afUXS9Vf7pHgsa3eJ8A27KExv6Gaw66P28avumx5mEA8lAr0DiPJ02
EiUF2PPVheNnEvAO/wr3O4ub2uqKBMj/sXdxCJpfrEtb+ahWaZ2cOe/dwfv7kPUQ
KIDNbpsr+syWu6PvEmA3WPT6ZR36f+1m1p1QAyB8FeDD/6/HjJFp6ufovZciKhKP
Fw9aDuNJpseJDH09aSIw1M88LA2P3MH6145dF/F2Q3+z6A1s9SfV0TJWsuILA4so
DklLVEP9hUNdNxiJj4zggrRpqtaMBPglh8yGKebHMVRTxo7a4qUG6xLDTDjpo9i9
CCblCsm1oi76BhcueTZboRXMJBN9ZzUhGf5ueqc00LfyT353C5KXB21KYpEXqFq2
jBuEJCRk0mM8lJw9K+1mg9GIbtBPnGSb5yb0ssnDMArc75xexWIeKHQC42oSHJ9n
gquwa5b91Tqa4ZPoTAyymnC+7kNsf7cjT/G+7lJyAoD2kS99qtELRVvBrmu6kHFj
D+lKBJklgFJQq2Lis8+2d0cNps7FYK85o5r8U4vEQ175+aNkJG1tECb92dam4TFS
vHyZ+qC7CYGrm0D67Gj8/uIQwahcMyr1HP96FwGZpuBK6kkVrf9+kkJ+nIf0gJnn
6EdnPcdvHBXRFjPTX30DixQeTz2qVzMZA2C2JGFgQdSBQa3QmN9w1cFKjbrCSfPB
lJK6fZUPasV7s8p8h+wI29oyEFO3mJIW6J8TCb5ION7/7Zfug6oPtLgeRHeG5spQ
3+3qfPWNP9syuj+yWgNsBP/+1ewKLGImnAA2gCXKib5Ddp2JsTHYzIZxtYItzWig
9+iit/ER6Gvp7xDpr8A93Tx0AUL1ihKjFkP96JF39ne78HLxYRiTidMXEF6JVRad
Hsa9zpsvUgJkBS73b4KRVojWEluQBiDxvNCV6SL/51XLSUX3HiEkXCHa5sG3cskX
cj+0LWGLHZiNKBrhI/irfNwrFWfud0bfgIi4fFNpokMd0jqqHQwMLU1mZ5gOpCDo
DRjzsY+Qt8mdlRDgLoVl2nLNYdCVJKQ+He48WpbLp8w2IN/49BaKrs5pARCTIDWA
EcQba+MdolJuqFXlPfbemK3rlmbV4eGz+UhyrCc9y+MYtG3PaC0PqjIWmGX02I6a
kETE0btkH01RlmVX9NW0BO77ZAhc3lF4rMfZgQHJPmoIrTbD1AQ2jvFYJxbLZU8O
f9DqWO0fJFTovgIJxPkebhYzBSItLsHr0iYewbjcke32EDjIhDJUoRilqbFTZlNA
78LxGG6k5X/7cMuscMR0oIsDN0QQdngyg62Z17oNT5sX8ve1ameSM4YmddybwOsV
eDyh0VAD8DlbA5kQ7/psmA+m2re3uHmUuLMeiXcKB2sFET1hoR6GL8bH6avfuPTV
nj1fLZHoB8C+6pXiQgsEyyHT0NJlIzejNXaX6vYn2FwKhcrf4kTaH5T1c3yrpc5U
AV0iSO5fA8kfMc/3FBXEzy5uIJQq0OgIQIR/VtpB6IHVfgVziIkfnHdI+/iGUwyx
XL+qHwPd6/uLyw6jygb95j70ePiDda9lc+5pGDUU7gcUhcUAEFZKy/geIuzxg3EP
6IFGH/PD48w4DVhISRYPhFYjtQeWdFmeSovKQWV52VbIDRwLdDrooC+kwxTrwTrr
gkaU7ERwSYxiJmB9CrdxOsHByFCXJHllTDyKcdC9/87shj+qx1tZPnnUHeYrPFBe
wUsBxFc5TjP5nwKwBOHyhVNHMq2NuEz9j0rEg0HLbrT0HGcvpmyJ1mlY+Nya9yYo
hcJ1V8OfCmV2fVtxBvY6OWZzF7gOiVDcrgvhUWsHHPccWZ2fwclsYnK/FYXv1Gmx
3A6MIXyUTOZPM3zyYHeK8KH5oFhxEJ0KCVWlFn2zQN2q0Mtpseq4tY7fwEpmfJvT
UqZ8FEUPqyxPBeJOeruR2jX3bc6Z0JD3gJDA+QaG23WgEnNMsK4fdGdiSFNWXdI4
fVnzw5AtCLxi2vm2hbwAB9+oDyM+aS6xHFiGE2h2FQUWfvicdf9Hhp7Rn1iFpCgK
rFxADYoZQPm/THn1MnMsYYcy7ZDCADMMnfjVls81G3VsdancTmZsOZPHj90mf3r+
oUDxLC0EvByGCCg74qFS5QIxUG0KI4ETCJSMww/0zyiUt8RMWnySI/8fhEKUhVF5
gWe8auNIhwptruzxx2fSDXLuyPvuYcvhp3RM1B4EiB4LEEcmmphEDfCuUDI5nqih
5c/o75NspGcLMtOyUITqUNvzkUQNp+3+EhcjdQCt4DffchweEXFmGHLWSiRqxDya
ATRVJBhzUeppYi288HdSqCbhCPEoN8r8B+pJZ7lWDrAYZ5sc06lh05gHm/iT/93O
YdGgIPRdWGWhXh+8IxpTUfHOL0WRkfcQIxyLUUGVMRoKX/z6afo2QQRHZ23ohuR+
WNplrIYHX9mgmTgYv2tO3EeyL4GYiEp8DXjTg5+JvX6Ntk/JA1YCyzCVFlYngnjF
/+trjOrygL9yL+jpEmbXBARVXhYPM+4GVVdukNk5v3478u9ZOs2T0eR3nE2XCQlo
T+st3pp/crCHfacUPr2mll+Ov/hOAgCP/FN+zVAY35um5BK0YfFqqq+AueY4BsSa
st/Xm+FIv2zkG6lPvVhxy4LRNn+dB7sLlZFAeza/kii9fjx5Nz6js0fMGaMjyEkv
SMpp7sOIwZGrVBjTdgegcpBvC7U6qqKC3sVvaoC5ygOQoe/p+3TvxJnOEIJYnQuB
Ic7ogoChJjz+JG/rbpU4RdGdmxI9SEqWff9uktVXPfNqc50sUwwkzHIBx6AN9W7i
HCoP/i5qXlrfhiminFgdwnSmaOWnMAsSqq3Px1wWJFC5ch9Z+8evEW4KXnWe/dJ/
Ev29y70+rtXQhf1n325RtV6H4QcnQHRAtBCFmf9D9DHf0rJr3Ye9BzRwgnkzETkH
9I5W8zEfa96PCvLtFwii3FyZ2IOmN+Yh4PDyV6A8kr0iAlkysK56lpycbJasSyd6
Rc+wKv4gDk3mdme2VJ+fIYsBLASa2ijTa6Yx1GrtD58+rvnTEY3k93boErmRywTb
d7ogReyjzvAfPkcGmgMaZ2UtWPfCg4nlDJjoZJCYlPxvTDSixtels6rasjhovWnP
9O3LFHArkD1ZiE3v1i8bvLFu7f2SOr7sbOl2QL5u7s8Fpw0BQxgVd3KDkOEwjqGN
5KTwJsoGUyW6pg+UCYjidc+2ikLUdxJLJcpy/F8OplqmzhAOnssPjnDfkOx6gF5a
Mx5kWnKQGRIlV7WMNz6Yj0qMjUc6fDcXabHjr6E759OIXE8bWPpWsZg0cc51uMJ0
tByDmnxwuROwKdDbWcWtQonlEOoPUZy9epyYooEvwGQ4kT40Cics5YD6MWl+TNPP
/aVsgSzxe0Qdw6XKgYh33oLF0s9A2MSs1iroKGFkp3vD8/Lkom++7xUUaRMT9WOs
ut/K6eeYvneiWBTK4t6SD0GzpixdUT20/QYxSNs3mLz3VLbBsQclmNuXp/ULbYbc
asFgD+B4aeAkBXwyc5FaaI6VC7IF7+JZRjlm5hsPfc5+36XoxGZpSUcqNzJPhdg1
ccasPW22onKiU73d+85gnpQ1TLWfrUMjmfHYTyC6Bb7ATyCmTvHIUYrjPy9dJLDX
tEcIukp7lWD/Gc6EpppzaHJDktTh3SuubkhRbUlcVJwqq331whUA+Yj75WGcOhws
rUFBD7Az3M40BnBvwlRRfKDmW8PrZ53uh0Sunxn1kTqhXMEl6q0GZGRvmCX5/FmN
M5zJT0dpI/duci7hlpdXZKjBQSLvEp2+JVGdrozh4mHTIPlXH21DdX3SzIRE9iNE
CxpXwAsuEWC06UPftNk+X+zFBchO1fk6dHoOjkH16SE7kiVJv9hRCcfMZYM/QhKe
/gaUkeqgZO55lPDh2JCKUczO9ZW8ZlS4W78LY6cDQ3Pb3qPTMiY4csM4laVkskNH
j6SPcgHULI2oVd3TbKRjK2lgueL6F9xWNbWuTPzn+k21P62UnYpzZSeYnsOT0w8I
4AdcDTjv2xOMzR0K6DV+m3bWljvXJ3IVFaZxIRIfNxs63GW8pRJUiHkDQP18HYp2
9ygVLbuyhdQYA7O+aQ7Z29RvCmrjmfS47TQpuzFJEUu1UjVklP9/vL0lBTgPM6yr
BbZSZGBg29MunPhIhoWsskqxe8APXapYH8WDOZGX1f7P78s8ZiKgIh7m+QAYLMg+
eSRBdaEuI407TKiXyH0MBlplVPXRb3Td+KrTOhkHn4mvsWCTyk+XuvVx2oPxCFor
iCilIbtLuV/u5XMEtTM8Wz5J2SO/vU0JYvCTJPAHBeu9u9Kba1ajP8zpVCzzEOns
P+AIydtrwYcLmMCo3pZHG5hbSUNpQey4dbQlKj9vZyx2Z2X9PRVSPThN9mYj/ho6
HNXkqu1W+yJE0P7zHj9hu0E3kOQk2MdLP+Bg4kbUrCp+LBtvhcFgvVbGT5p1KwNh
u7UL7Ik9rymEWT5d9crZsucHfsodvtioKYqmCtQpSYTY0nx3+1UJmjKEPs8pRVu1
HtrWSP+vCL4OVFA/gLicyNe6Z1hevrbya3m1QAmy1bIQlh0ZvPnu/PnifS8d1vCU
6ngSnCIhQP7+VEwB9HBbLQE4zvtKWx/58dhhPoGRXWWwl0Xq5K0XV9L32kK3DiI9
a50EgeAXvSl9uF4egn9VwJxP+3Abvg/vexE5OdPb3u4Rq0fk8eW19qNo4Kx2F0ba
VNJS00Dny+EwcWgEbhglP+HcRy4w5q6R4pJrByWp35ivuuVO9PHik1Uis+EWVYRe
C51QLyuyoGArdWB9QrIVlntSIHdPLgYMTw8kBRdkxxlRfx3Wi8Jh/wv4Hr2NdmvD
TfgsWogN+uSiiZrw/jliMiuqEFsfNNJZ1coBganalyeGHnmXKWaHC3j5ymoIolQg
GE+p0gOT+l9MC+C5Jr0L7Vae7jZUL6Df628Hlxsq+enO0eswwsv3UJiOUZ0CCwZq
Hr/rgEe9i/TmWUXbGFsu84HDO8TKAwuVJdT09aCyxlMk4mhhor28kIdDQR/Cq0HB
wNjiBcqzRO0QGj63P0xjuL58o2M4THmhVcDE8jliRgwcDFvb5kMW+s5jTs4ko2TE
UpG7XpYcjpLBNZK+thw9rxiEmHGNRmY6E0HRZ+k73Y29pEA/WSjvpYyU/y0Z+B77
gYiBquTm/Vr81XZRnyvkeIsHPeUA4Al3iqYQ7xtt31V2Ef4xmj5KCOTBQElNOh+v
LTW8W/DSTYd0wrZAbEMdaRBrXR21sK6I3RmabsxEZxvSu3FuxeqmBqCvMFLo1tYO
IXyo6WnWMEvRO+5hGDbLtbVFwerCvti1vrAd3Aw1+gKsormxrUHg/pQ65znSyBDB
aznV2OJ1TzeW6XUwVC+1G7C2V31OfSgHr3DvKbC4GV4rw3S+y/W3Pu6fpyACQShN
bWUkQop6hifJNIx0IK2yf64o8GYzDK21638Yhy4K7+fLQdO5ftZnSTROXa27ik9L
CLkZz46cJfRyxhtCgJhF2yWzLX2XHc7Q/KoO0URhB/N9krN2Y1CxjOAukVLCmMbZ
/WCqLbPb/xzXVEIXF1vpc5OjCTcVtGtLvPu/gPfnALxmbXZGP55OzEmYFSgwfWj8
SYCOIht87NXKxhjIJKa0/ksUyWU2CoGjMMD37N5obXLbJSep39m3Ak9RqIs4njq4
0TWlMji5gBAqSeAsH28Qm/RgYZWinDA1FYjpT5fbYusn7xZ5vtmlVKObg7FqRt/Q
Xr1LPob+w0tOmXuCxoy4KmVVmmBm9cRJxyVrCjhrNxLosKY6wV2Iro9EU9XmVEOj
qHos6VJWW9q+9wy5nBC0+94UUI7iHwmTcTiwTDmdHfEhn/Es/t+Rc63avyJg9b4Z
6BYnFVmWHNmZjSuaVJ060a3rpW2z8zid1/dhO1Ww7Nh6WPk8/FB9swZazZL4rMVJ
aAVqIJ7yHaj8aCb+3r3mvDyiYeur6wxj7eLoeBOAbXcnRzE0HbIOK9VHnDycqfOK
hEf3UYbtce/y7e4Och6TZ0AXyWhx3svr75bqxIS+pRYYaCZMB8C/StaR1AOa/vdR
hq8OMnu7AA8ahMbfrY5jJiEDcaK98gNijPttFYsezew1sdbzJVAlKB9z/qCxjgZk
O4hb88UesbiK89mTFiz/dq31raYwtdk6Zrhy8km6DOMGOTr4Sgpue9PYeUuyUYyu
YJlYl/7MtW00sySaPtzUZNEuKkCrYO10U0AQ10g8C5kgprXK+6DkspChyeOSfgpl
/1f5FWqHp8lQ5nG2W6m1QXPRaqXf42K3fUANT4XDhCmYsqBHFXZgr7roOaeCMv95
v3xdn1Tg/vSFVorb9n+66w==
`protect END_PROTECTED