-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
q9DlumNOvWb/qgYdd+oJBtv7sZ+Gk9FVhKG+bUxkERZcWCPt+qUHiamHpSvXmnDnSg5sLOzgIJ+y
okVKnkGbtr1UAYQQs4EDNnRCzKoOq+eIcGedu4Twj59CAQgBLoVr233W6fwd3aLw7p+fsqRY4NWv
5KUWJe6bU9Optl1zSC6Kzm0pndZJ8ChJlfz5C/atkq2OT2qF2EUB13aFvh7P1mlR4xwrJ1c+e58H
+mcdnI7AUVKpFz5xvvF1+d3VThsJtlwcwxNSM2Mh/PKeIN9qqDz8uJCeMulciLGXV9sfvuAl6cTH
bRafFhu2gMYjdfaPAbBBERXGFRcrOKLV/+oOAw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7808)
`protect data_block
tSR801Wb2OBIkcVyRUznAkbVVbmYKZ+m7XrYmpxYEx7252QtYFbGxGiWtNiM6w0Voav1Yb7n0daj
HY9R3BSCBTOwPzAXxSJxZ7HeBmfBNlcZ5+w7DcYJNzv/NXp3sqv6dxQMP/CKbK0765uS33wKSUk7
WuNBsTpk8qkM+N0cR+0U45heo6hR+cm+YNQo7Asc5hthZcYs6NtaL9BQLpXAIB3tI/aRW9/E4XqP
NKYscv7UHM3kZIbrTVt//XMlAKJDB9WeUtii4Da7eWXWFSNQhc6RezLPGAcoz4WYYFGfgxKy2mt8
qTypCWs+jj5gM4iG55JOVYNlF7l+7w+/+TLY4r4kdGP5pWmFYLFhi/eucArfaWpHlUd6s8R/eA5L
Ux5H+dGqHIKBNuA+4/jkH7l3uqADi7SXLCABOf7pHDvIWT7BhxX5fK2po0/EXH71A3f3/MmJvmJz
sscLGc0qp1reogVQKzuOW8QHCSpsqXSXozpCcIIkfts5NiNpHB5TgNmDEW4At2KX/++jwSsPxAdV
mwnLGqyEeY3+JUSFkeIV0GRFPAI4Tb7PZhyyvLxSa7QUTcfn0sBg6ama7nb0TH/2z22SMKElApo0
eF00AOlhgk/EvtPOuapTEbycFlP0wxyiALX/H0juDGUEDSAf7HcjXnsMdPmrgeBby1ncGHrFzp+L
1cqPFgL4p7eDhENVRdG3fia2eMnd1dnHLooyIVPZSFk409M5m1Q9T1robAJEwf0wQuE0dyg3Q1O3
22AvyVqnoxudwiJ7RYfqGF+uUHffQagiJM9SqGnkG06+wmVUnaooiABtZc/Y6vq5tqRezpdArJoz
knY0NxdaOEfDwRECIYr6zrOwGFwnrjNbH32ThgotAhLowKG7updANPN/3hn5XcGD4mCccoWredpM
mRLRKb7HsQ5dRtJEgRxHGub5MT8GD8s2wAiXshH5t1gHh0bc0XIJLgU9TR83TiAbQTPY9gSot5uo
AcN027y799RYetN8/eh/vuRMjhD3dikhX9XzQr3s2rhccsMemvxJ6cwntztpKmXg4PrBUUYYKn71
0uAm/TlihWKnth9mwHItQX9EwWjGM8/pLDMb1jDvxbHGkbANTpTY2BXGhQXRCVesuV+90SezSuLu
QKEsvme9rRftO7rZNJFXV5fJ7eih5XfWtvByqk2iYlKnQbHwn3OGe3m17+9X1wX+lHHcQBky1tjH
C2hLkTlUBZ3gc6mQNaEf40KzVwf/TdIrsx8FwP/hTFLODdVQiKocOqFnPPIplehYRgxmialDRL3u
2TqAjofOTZ7R0nXQW/RHjIdzaYIcygZETeWfMdlbAgvnx2oNP1M868SdxsonQaHV5Aq/0YJ9Knpj
5XyN/1JuTNNZOJtLL+2M3NXg5k4qEqNvMye9Q6DqtC/3pyCb0i7mycdkh0XZaOHK5Neq7u5yd47m
2Y+yGn+FJOES44ePpOcyit9C0bU26WN3kXD+dy5/QxxvxqfldaX0DwcDPtv3OsDIf8H6PPdfJDz+
wPUDTidQbgWf9Fs8mmx1QSq2M2spyhqiEh6IdQo9I7QlXg1QeK9/YHTrSZ8rA5jyGYlVZsN2hVzi
W9c5rfuZ0G+/8DyhA7P+DF31gQCXPS5WY586FDrERzNfgtWnY8Nvc4GN/a6Pb00q4jXEXO8itqSz
MmiZ9yFa9xEDnO18LJMhBfMtZ/nocXn1B/Vbv4uXTaPjVPuo2No7ib4PAoprxXsb32XXZhsNiveD
0NsepY/FgyD643BOeObDN3tZstX4S9H12gSeYfiBM+igxzN0tbsqbUydOb3IAXDUms7IZbdwCfCB
+klmznHeOLIX0R1foCqvCzFhjFmoZjGgsxxcg0NFaPYXionIudfaw9LNRhMXwrzUc6d9mxkNju8Y
S6GJOxJuFtjLQ2fhs+oO1w21YFWkhhlq/ccpKSqBMwiXGRXCgCYlrca4TT9hyZgkMHQh8ZUWcQUP
j1h7xBmhkDuTVrsu3Evr8DJVVRsgIrxvthEMy2Ix8bqrPGLTx0q0yTf4yXDGQ+ilB3VTkw3wF9Gl
oXSwZsV0SshjPQLWyjpcGpWGfZ4znIkFWaanCAxMoqV6mUl1KBpKSoJClpXoGlyH0DzwADl2kuHE
8v+KRjPczNWIKFECwNK2p+K6ca0/66U1jK2KAISjc3r7pnySxRuryLEZ1/mNU2nD3Rj4nBVY/zjt
yeBxx37rw/49zGmPun2FRNfN/6JH6WCv4nZN3LXuoISJZRRUG5egCqub8bn20vPCNp8M/6eYVMf6
YSYbKT0vQelcY60U6SSS5yr70/dVRj3ZLHJud1d8WEIpEzDcKZdhaEdEvbK4b3yKwlAGJxX+ogQK
OdfLT5HthMVMB9S5un0ECKG1KOkq3oqNse75QXidYdnYvP7vGK1AP9/f/BVqG3AJZoQFGF0sImRj
7iOrUSY3jz9NhdkLZufmVRpwIwc3QLmHnGKAVESF0KYYNj8SjVITYb50ZhMYxKKA7D0uPq/dzYCh
sEQTE/DLCUojzmsjSFPi2UrmE3JZTxfjz1W17vATrEiHS0UhuvKVY8Vhhm1C3d5MJMrYs1f4Dd6T
a0cnQlYp37ucSBJuZbpRo+FA9JDXgEWpsWr1DNSyxY4MnePMvhNVBtPL3x/Zsdk+vZe+R5Ldwiwp
yIXdWHUSgKrJynGCJ/TAsjziXqi/0UAwrKHzd1IrE8WCdqSY1AK/A9SODIY6ajLIxgEg0tZaynE/
XooDVxPVa53/yjUlNFWOJbsvnSJtszVtYveKd+Xw1btiIQGcp+swBDrM4Z0U6LQWXCOjA5pBDy+8
xlzPW3UyYPaIauCZYMF8LGfEVYlommLibxug3ETRx+Lu6Rj83XIpYcFFQiPvdijDOC2z2ZXO5cak
lAGMR0NdG/5m70GQDLJqVZHg7XJUMeRAjb0wI1f1bkwL4MQSc3PyWjPpvtmhvSXNJMXmKytP4m5k
pM3EkBrEilAdUpCdMUL/WOvNANCA0h2XEYzGsmoi41Y3o+ih3biNf4hByJKHuTS/9H1Pzyk9Wtg0
nQjlgtgvFoSSXxAV0XDxVMWJ1cxeRj/IXiDduJ1ZOdaUQbpsV7C0yjsjBBfyRggFgnDVSlvDpxXD
ECTZZNTQ4Vsy6kybUQiaW7paSbyS+TLwgmxQiNYafrqgUezl/eWmg5XirE+RTJXyJyhupSQwu3Jj
8XkN4gl1Zy8YlcraTdoXZvDVL7VsaDXbqpKnlowNTKKGliAgBVI246kcOd9MktJRZJZ4bGehvh32
FmWItCC3cTpnpylJ+dj4im447WNNp/pTeQA11n5uxPoK1mnsO/mTnHz9TdtC2f7344L+YpIbMv3R
dFVrc30x+g9REjZLs9s1H43xSwSwY83gkD1dW0M5zPKmBBO1YfWBow45o/unLNAL3MSvMtcrwBzQ
xUl58xDJlonUEgucHTG2HKK18C4RiRXTrA2evTEzL+6lQO7z5GYxpvXzrA2IpyS4eO3oHZp0VRhi
W1J9dZ/NG6Yp18pmF4gqpy8wOXVZGt2RKsOLjG3/j4Q2ikwMpM6kJe5rQEHc3JTYUt9rdnfbt37p
wzV3EFY/2itvduQGf0R7Qko00Agud7ZsisqAHjTXT1n/FpTo5tr0fXFIvQyBxqAbPqmcrXX10mIH
Js3LaWR0k2haQ3Wz04EnU63KeFYsYdGzlqPGB0A/qrFHbvVRbTkhVWedtv0xknO0+p5WGEJOb2on
qO0pzRGlP5nI5+XNEy1ncvUvRNBSF4CCPGTLVF4Lif2R3xfMB82OKfQEiKs9C0vyN9EpkdK0L3h3
SRah9UfF10GFlnN1ZgiTRgE+/VF2oTvz3XRGlF9Eo4v7I8p1sSodlxl+nWUhGTMk5zIQlmY5tOfc
NvsEeCZ4JomdcqQafGBeKqYeSWBUGizNMhjAOGsOeHj/DIHajXZaPysAKJg3/tjr1gvH/3C/QYBm
pZgySsdcMhAdcKVxFTEg/ydUWSuEozHPIjhrmeZ+wymea53+FkGkmOQuuW1uiC0p6OF6GrTZ5Av7
gVtky97DkO1U/tlng6goOpDLdaInMN2HJpAWDu9Ni8z67qyKUkxeKL7aFlVoE1vcZiDWndwKwqUy
eqO9lL1In06G111b0T70vf8jgtW1Egjd9A/CAwbi2ayeAtOZcxJER1v6YYbWJ3jUCoBpb96Isg64
f+Ck6Xmya4JP1N3bGnmFeMUpbD7ftUPqib7mIxb0PXYClTnexuYBsDL4AYGxN83wiB31blEZcFf5
a2GM5IDchxQnORtpvI2UZ0XZL/8mlZU/He+VcewZaBw/y5tTB+jwzFurlxP+gbUlaIv4icKZLrU/
6VLGxuD1YWbBIRSYJS60agpCg7lT0Dav+h2RMkseZzCBfWzoGPIhiGPr4mJ7Bd7QNt0Ejfo956w8
wOLKvQesWKpU5Zr8LjV5AnY3zoPa2O7P4esOorzyW9a0x+H7u3jckpc2pNlDsM4tCl779KrZetOp
C70Jo0pupkx+CavQLPPWEtgIX4+ZgaHfuiiVMok/MJtNU7xmGPcRihwQXLysVAJAf6S3TfsIFNft
tZQUtEE66fzPqkQbhRMkN7f4S4ydL3avJwvo8p2cVszV88EFb0a60qxAGEIH1KpHL7rRD5ebNCYN
q22sMTr/HH+A0wzd0bKI1PJaVkgxaTafeLgUKfc3+YAhpe5wc/LLeJgOMbS5a4vIWwsns0wJLq08
0aT5BEMNTYUNY/T48m0y1PTbkElYHqJwY+bm+TnVHwlckpJqA+ApVzK9WiGOqYb9pRwuMhuO0RiL
1qM7HZI0waKsKQq/OfDuqfOqrJxYhsSUPue8bE4GA3Op3CRLlS6iVuUAGe8CGGsl8+IMeIALKQvf
PxGcSoW/dIEiTxStTuIRmmLWn0m4y/zJw+Pbz3LZr5ypSHvI4xLtd8jRjbGx0YbgQnJAthp1nqtJ
5mVwJ94naakmg5GBMuC+zlmZjW11nbtG01fiaczM1q71iqCPQf568qMCY7PVPnVQ5gq516pvEcTF
S3lFBlTYbvZ68xesRVrKOM6daZPe8fsSIWWwqJ0Yk5Ffr5p042EFN+TiZE6D2X3p7HjQUh5lK0bK
B3yd9Q+RVmTe7bUG1YZVuJaMENDkSmEeSIN/mCLieB5ZnwIqRnWXfmgYS56Tjh4eP1lLYM0fIk/a
HtZE0z258N11E4Wm/QVwBW+9KvUn8Ft8D+Dj3/3mzw1naL7jKmumhkAkewzZXio0SPoqdM7gxLNn
LKjSt9fHhFHlkiP+Tj4oUDJsQv6eNBKP6Ib05/4BjQfVfiCdOkuAbt5zRGo5fVgkPQrG5x0JRLEa
A335I4fIMruuDBfKF+Q2XoHJfBmiWBa7gNkuT+6HolHRYndybhZOdqmv0bsgFNEQJwRiP+KxR39X
5DTzqNkzWvwavddC0RCIA4OEF3U7FLLITkNysqiTpqfTJplKpj6ql3hmAIBnsLKy5/Te0wWSZvdR
jk6oIPBR0HDkk5kNTrLJ2kw9NVDdj6P0pDuFjT58x7yH5cifn+YUPkOuMAXG41p9NYI8D4dYu7qP
4DMiDy38cuWy6Ni7Pfe+iVrsf+ilSb4acHMQTLaTVmsPA3EiwQVuyRwfbMNIDU+Tit6AqzlorxdC
cBbm6OSe2WctOh/4VTlpeOEOmoEveKFQvshz5cZfopTD+GJ10ib6AQ3/IHX7v5pYzvqeoaJTWq56
4L7Plg2zROhJanIwbpJ9h59WXZfR8PWRpRaVWTTHyK+Clf3v4jpz8QAmg6mK85jXWe2hPvaUcjD2
W3oKcXFJjnRWPwMn8hB/gIa65c839UoZloNdcQv0RnUtiLGeiJLryMq8d5w8X53fscly9POesUga
ZBNPB0ifXVKb63M4gNHtsXOBOB/ePI/GX7h7eYZHYFIaQPUTy6FxKA+DpDt0x9cKuhdbJD42fDsD
LQJ3BRd5iSrnf9h8oFb01CzJADgaNVDNzMlJQzOz8nkowgnqwFbN1S1N064ASEAIIAp6c7Uo5h+u
P0xPViUXwVZDWqgNusmD0PwtazeMegeerRDJxiiDDOl+AeK9vNNzgWBZ+7qq1VrRwzmzpII09ivl
FPijjYLWE2k+m8PB2wsxHqVY8Tj0WcpewiTVLADdU8soQPeE4okcm4sXeKZOW9PrlynQZMSP3hj0
waJhWmv9BiPzWvL+gE87pkQTvuSh89JXducUqTaeWTTCQhRmKMn42lNvUQcswUUJDH1bItAmkA6V
lB7hWCKYDGWvBIlXY7HHZ8fFVjAMFteaAkn8NT41VIEbyuyW1XHksYXn9fldv9uxWFsG0d+01lza
3ORLZF8oURhUA2xeOBpL6Vl2PD7TV0ckKf0MtNWHCfdVuNCK5ggdakYO/vhq066lgPVjdh9GGw6Z
IY3koEh5VF1Bpc1j53kPfqhL6zp/UcvIs/EjNyhH12QxVsA/QvoxAqp0ifYUY8+ZuKk/F71FCJkJ
NTmIdEfGohKiP6X1y8TFb0Ma8c9ks1oHi4MLDPDR7fCNiKAX45yU4ItyYp+YDeyLZwlxdcrwmOJU
c8QmgRZyyNJ9V1w9zZqxRJuPcp5gVHdCUqHlCwvoH67iNmEx8k9W3p1qszfAgWvh0EZB32hly2jg
TjFOr7biKrf7uYo0PsSnEteZtqQOLvj0E0+kscfwMTOegDqy4LGl1TieCa3R/XEuSdmWXVEZWDhn
CHAxX9lvIpxbee1kOo9utZild/u2f7oGcKq0niw2qL88rWeip1/3CsJG/DwCqmbFzN5+r/e2ekd1
tx4yg4GFk/DiJNO545yLGQAXRRV9Z/G2OOQguu4cFUG20jzYU7FVeB+Lb+bQvRMl2tdbzqm+WtIk
x+JBBmwgnb0hqgyk48Wf0KktTxyGnFatFMkqctjKCjg2k4E29osF+nwk5BCyEcmEIsF9/9uLO4Wl
DyF9arr9KSauCqd00ukG1/Zh6o4tuD+f4VoNgT9yUDKDhlRnIl0haILtNT6flsL/j81n+sX5kCzg
hcMk/97oBmz7IdUgT1v8bbKNRpkKinoXk+QHh9gPUm5CHfxAI6IXgt5ug4ecY/Brk3ClQ7s3qG0w
6/L3PeRy6Ibi3T8yvOO7xoLQvJ8mB+3M6oWPBRUvL5Wu2wgkZ3VM1b/wv6xeUoznRbBQtngmEn2A
nm0AmZBp8E7I0DXV19g0IfuXPmjh8cJvYGeyMnCibcOnApUv7lbWr28VyuA0ebf06oivcWg5Vnp3
DN9JzHnbyNq14fHADp/Ri/x1rQYWepuCN7jdFl4hHuNshhGVgm52lD3hWyig1eP0eg2lZ4qpzbN1
reCbSDrjuK/HzFPevBgJc5Tra7xLPgQZY1BlmEuVprk+wFGnIVUTn1j7r+CGeXMbfhj+1ksOXa9/
U9Ws6emktviutv4WqJETMogA6imyNGJrFqXVap4aczzfnry3pxRTMOTRRXL7WLhumsaSMZnQHoCy
/2HpEjcXS3SnsQMEAA1dPRbKN37f/PcjYyygsFP69CmrbfbK3hRzP8s9kGQjY0ofLj2dX22ogxNn
cfcQ47GSwDgN0BcSJ2IDnDX53B5Dc1Chevkep3ZDk/cES6Q4iR9vWAMXGOD7p+tFd0ywCcKQbN1a
N3Pq13urbz6UvST0Vr2EUBy0unVNCosKwtQZ0RPSFIKFRQWTXc9zEm8vYoKvAaRFFUZ37bTNYMaM
zn7r3xfVc8xCYaO9m4hKa9kjqQKIWYKUWWXB3MErxkdvPwix4KrjZMw3AC75TMuQOHm8MZ2zTVN4
K8R826OahT7TfdNu7fWKaE57SJqmnwBwgi8ZOUKt3vA1WL2KmFO0U0xyChB37gMpeBbiqSV9LDLx
TzSdE/x3pBHFf5wzrSVMwf7LJldKVRo8o9/ZhAO3wj5TnhMojJnfwBVFrb0kxZN7fi4hRc/Vv5ox
gPNC6tYN5QYXd2dFdLCWevJ7RwKV9AZJoDIma1zZ67H3DoDHkUkV/po5P/5P4qTbwN/eBSheIMnd
gXGMnXyxZyCvL/wtHrWOBSmi5VpEGsZBCpLUb3HPQDFzqlT8VT8tUAEdXInbOEL1qXRTb/uRVz2w
LwjRp81ojZhHdIzkOIkR1wHL3f7m7WEjAog8mGfL/G4c9wqiGbwleLHJ+JzzZay3rDALZ3j+QSO+
NvcIoRLJ4BGpxmpfP4MUvexqLcJfcHVMqa5dfznI3fcyLD8JUH8E1hc7VYSogt9PAhN/d67ntDWz
H3rPzSeQ9JeaW45bGXZz9rj2YujwWL6HPi3lsEWRuoBbRgnjiEvStpWsc5EBMNYs07XqeEn0qmC6
gPJ0PuPtu2UHBQr+xceWbBtc9MlTDP9CzVMCR0hv1z8RbjmpA6QrII1y8Qoagt/WaW1z2YGaE5Cb
behbWdfeqf3zwDORWrBL6qsRBnPXThydz+kI/hoF1Mdzsocxenq+cAd64VyjRZk1i+fdCA4RWXrO
RJpsPKGBb2yPqp+si1+eu5NthGHp+ZfrC6wW7F3fA6oN7AYWCT+lQsZbg9BF6knOWCfE1JdLN1tW
JGW+aODtxtzQhk1Nd0ICTWFXjB7dKiWRhgVNDOwcCJMarWiqXG6V9ZJE7WHClqiml8yfVbDhvzaQ
TZpTT2NK9/iHyqRYbIjmPTYCG35+U3nKv8lOtIXyUrEAqCIIZhhDyPo/h921ZvStehVzfCvqc69D
h4QYuoglZzF6bbquKzj1Hlc38y177L7mUZE5xCWbs59ZvrEYL2ZCsgvMUJx01eRGyhqRJUPM/2IG
f26UjnC/jLJNpmrcKWrJiZF45Kr11KGo3R9arWHb0Opb888BWV5kVXa3MgL0Jrr5fqEzBwXTdHlF
MdbCKD3ljaNtGWbXxg4zRl4/zMtAmiQqgqX7J+CoKJki/Ur7EGT4F1xQOILksW+vkGgU5ncKFtK5
ChN6guQgjkjvN1YMX5x+1FwncjWKXsrqoVJTVeS6ojVDzv6eb6h2lzskyp26RivKJzriOp8g0+nB
lzrMJLzFsSMDW0ZnE+bEjQyPS7ZFub85gCAYHrbwom8OvhdChLDr0oKcI4PqVXBfk2J2eSR2MosS
jM/rr9+SM6hU4StEcF4H14WXXxyhNyC/SlGsuoDcvc+/P6QZu6FlDteAqWTuviJS6H1M1/IorY+I
+JPX95Ja9ZppqL7VIw9CVdiWIWKXllytqJ2rAnvAULOZlbe6bPiMDEhavQwQklEBMNpWVKAmInPl
tUciWhP5lfWUnlytSBKMwfRF/re+AwfamFOyFwK2+y0qg0PhEMFk7KCeIN9se3wufTGMXvMsoB1Z
qoOMZmO0tOIfCA3X34IL29y4HCXyGbqq9TQ2f1g14nry+UqvsPvVNjHJTBazIiQAEag6OgiWntGd
tRPfESDoT9o+NdCAXAKtCrypOZv1R1y/QEjB+eNpRfEg+6ap1wSaPPPJENfhEdcB6GYTgucnARc7
IR1nkDpT0oSL5aGAY2IrZZyKoD/ZtN8RUyazXyBydqBcSyD4MMVGws4KywUuji436xOOeLByDBNk
pdxBy/umGWk07MW1zF7wYj4aUybhKQNH3+Vu0aDhRdT7dK20tQXcfk4HqKyVnJoV9LC061kgIvwC
AnT6M/2tSUJCicf8HrmWmlX0f4EDt+zRBBLu36f4E+jw76xDf0HbanUaO3gqAp4mp5MI1U9PE1UT
K4dCV+XtNg6O2LJrWziShHH15FhXv9lP2ZoCLs/rGoH1IlhNCZy+CEIo6j5g3cEsnYiHALt2yfdP
y2zWKijubvI//TF26O5BUPuzIR4t1ym9A8zhHfPBG6zcrFf6YARIUbhZT76xV6L1XKE+cSDgOk5k
ASgHrPQuwFFS4WS/2MgIlLZWpHk4KHzo00zRHgBOa7Q69tVJGyvEGX8Gpodu28K11R9fG43tKP3o
J5xi39I0gC8Pxuenrqw/nOYlqNUZcyA6URaETk0DPpNxjrFkyjyQ58BVPv/erWWzYYAfxS8Pyozb
ChXI3HHJvWwjS28/Gu1Ko4ZL6p7R53D5dpptqSc9usSKa41TYAM8t6yYjoYzJ1NQJFmj7rmCi+jX
DpAVrIVP2AxOAqlg2pkiQ7tMO0g6q43XYaoMnqlhwBHMz5zVfRkdVLax+o1YGJAuoyBH8s5kScsd
sE3hX3N37uJ2xNY8h5AJesS9znVCBQmmFo7IqnlZsMpOjfHiTq9xa7l43XF7KfstQmwe+k++yXJc
VdN8JKgeKxPiCjwNu645SofdKHWLaS0TBgfcJnJ9zY/NItINDjBcXRVUj0zynnddUaOdiP1sU7HW
Ql0GI4SHVyKS2v3RURIaZDX7Bltoof38xWL2RAukOvI0XNjHpGAHjrCBj4tnUK/AMMsVAMrqXDKZ
AYYaszcUm83vA7zvNUGnCnjLa1vS8q0WsE6q/MYa5kvxXR8BwhwXhOhFN3yUjfd7FzZZgWNf4gs=
`protect end_protected
