// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Sun Sep 22 20:49:28 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
R8tHuOysSvQDwXV8kP8mzTCy+gB2pNBvLkFJ3angHqZ1bdy99ZJtAeFBYFjKletz
0FZTl5C0M36MVvppZ7EKnReXG1K6ZojI6Bllv8RhSYnH3+gotQMbm4Wlra5EiPIJ
ywJZewghf7/s1ZzEpMwtIiD7YoJNy2q4FgcswconRw4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2016)
P2oHQtd0m0ua8E5puwayd8iT+wuBe5c2LxLGvrrc7PjAGXMzO1bqqekTgxzD1mKP
5SWMaHH9I+4SCOvLqdUkB/0wWqmX5AQZwGJ7TaW7q3szuVx9w3krQkgBjkBb04tr
cLU2TchtyJpTGNFHbASdl1ogao1xf04SW2S8lslRXLUlWTNQUyJ9dVKgZeUt68jH
cnrlVkGGmRnnbFLDuUZU4U6ZQq7Ujb+lPakfQVKN0MdMHaGz4IRFIaH2I909Dgya
TdyDeckUWko2bd9J6ypBlWwHHFCgQLKcc6r7na6oOztpjulFgmNfJ7XbozbzZzDE
B60OV6G3wo+bjPw2I+193Fu9nve4u8gAQTBG2TU/8i66S/x5wdLkY0ZP+MCW2PTg
Xi9r3zML4d9LtASdsttqA0yQ6J50qkDqLihKXeM9m7HEWOYDHs9bKHwIY0aEPbCo
0PFJom+9/eHOp9ozhkuoYaCvZ4Y52EaYO5IY4znhF3lj916TfWW9c2IvHVTAk8kH
MWny7hCk3wkqf3BogPy+xePq8MEc5tA1dFuJUvy+WKlcxD8Zv0k2fV2bFEKFGMNL
eNV7po6DpJtcagIdrWnjXirB/y6h0GS3154L98jKetIiKNTelreCKypw9CuU5imf
Kbf6q0u/sO9EUUSn4tNDKB0hhZR8yS+HHEdAIojXsHspUGoHQ5Cdtbayq3y+dRYi
Io7MoORT0Rro7iPHgeBohkFzSZ060RADR2G5HsD5bA6gDJxDrrpOq1Bbv7UFQmpD
XyLDjyZiK/gmvDPp8qr1UOfU8NK0uMzWHwEX2PnjpVHsdT8xMYAJDO/ADAigYppT
EIDs1dQ5C7Ll8aBXYnCm0/mM67XCLly/NXGTV8K42yvOdaayjxAmyLwxcNl2iHIy
bT0V1596e74BCTpCE59K8pc02pcz+UIwxXfLb6VDl1RuWb7DpVHVxsRrx3tDR5JP
LVjodEjvhdDPp/IW37nqCGhEQpLjrOe7HTnToVj9F4BEjEfC8oNrHY+Ugdoja1aN
LluV7LHbTS2QFlXpUoI5spUprc7DitIR7tibhOqRNkbjOFyoTmbSMYyzlBjW8mNt
qv/RhAKB/MhEpPJ/MD+lRBQ5cdP9ZqrMUdMrj/yPrt0JVzewqY+Dv1nKrO/KOQ7t
5kFqMU8vEpxd6CZ1igT3fcrkZj9g89DpOoaAJsAuYHSVRLakFvyxwW/gOOXoDaja
J7E65WkfOWd7e14REKrq6L5wmFoTehhntflT5egIfw19K8HQsm+rOpAz2lq5ACza
A8kIuDKBXTIyE9lrjDhcyo+S9xtGx66ySqaHIT0UTgJBSzBPiwtp7m2w8BQGX2+J
t2s8rrawvgANezVDCT3759x92nZIK9QTGXDlq0ibOJPqc04fa5z8RPwvZ45VmbTT
RcgfnAymvbr/w1SFD30BaNP47vyLrA9/eE9QUpFPzM3DfycF8nljmUCVZyacrxpO
cyEhLtiSjFoeJAzXU6xLPaYc0eH+jo9xLeF982Afch6wCrDJJwyCwryTF2Pn1Rjh
Y88hESaT/ZFXENyho3laOLEOGSNQ+RyG9ajwEJOCt1Io0x/KncUv8R2cMLNB64Sa
XgOkylb51sMlHipNEVxnZgk5FCFGwZ8VKFTgpOkWS/IV7NaBxg/MDF+R/V4/43mJ
qdX7CGIg0ITbJvDe0qfGRfN7XL4BYBvcMpdWdDhb3qFsFt5c7QxQESqZj9sI00k0
Z8+5z+YmfDionZDLcdhVdLDfW5g/R5PS8KGdtr7i9jX2GxWwCFW57pUzUGrUg0mv
Qqhjm96R1EEXFrR7ptxUmPb7yIXC9RAbxk7sxgUxD6mSJseWNPHMRgdkGll6Xokl
mqWFQJTmTkPVENGHgwYdOOr0L5nStFC2EEinm8anSeZVoU/h+GuuAVLhe1wmJOYn
R2WJxdZk4NatPVfG3HaOYQBnKGx0ksvXZeZXiWh8x1QvShPwU5XPBYONTWpgUrEA
+Hx/z/QVrdMNM+UjdYwqEXroiszXZbpwANoqKjIxQkBkPzljtD7IwNnw+FdH2L07
xgKGsux6aO0JrEhwb26oE8xRO1axAlzC4Um2eAngSQwwcNYzq7e46peqZzpadeqO
gFIwlvDwIN8TXuuXZTDUT8q5gy3OOvPXMV7KSBsVlbUxWvRN0FLjRUmQDn3zFvx8
KL/lon9+282nW3nLZaADR+/iIt6B2EVGifdcNiwHqqieYNnNGa2iPonrffqxtj1R
Fgk6RU6vgRmzMYEli81qeNT1RZzYMXLWJ/j9Dl06Cb9osSKO7eRIYEy1xwBUhUWA
OAuJ1f8yukPXS+XjPQpXWe5WLfY03iDMgefw9e7VVbIEEDIfG13VCO/9jFahHjzY
l5g3bjBMaq8adSEgcn0OYoCaLz0Nzv/9mLTxSml4T0GeUqNY7onBzVc+nopuEowk
7rj6uIf0WQcMBN0ZoT+QYyKm/WvLwGgwd1zZEDz1YiVE9AEHC4gRvlOL4phpJOin
cEZ//AT4Pu7vSAhpbJqvCGY/4woaNLEKkdxu3zJM/M6bDX3uVztZXNy7YzpmYlDQ
XypQaQgzfRhHPF2oCzDrvOqeyBBNzXqMnYr9kCGC9Pn6m/XlHyTOb2tiAJaFcJdv
E6xIVlFIe+FW/ubvyRdwPx/glwczp4cqsTackLpGlmXDX0i7IXoIHchO2n44NhFz
`pragma protect end_protected
