// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
gyqwK24cmHEXPGhgUCKk5M0Z90iAMvJsWhwW2xTeQKbtFgrpI6hVdeIsRTVsXkjw
aGXvyPZX6xsqavdtae82f9SAwXZN2Vb2TMug8wP2mSxbG1P3teCMgVMK/YUspjwl
7pCI1GiWvHWY265z9Za3y1gH1g6NIEeY+YjUItzZAmUGmFyfHdu5VA==
//pragma protect end_key_block
//pragma protect digest_block
TqMs2cusTzT6IjaO++jVeFm7jMg=
//pragma protect end_digest_block
//pragma protect data_block
Bs4gsRmVrAFl21Ffg+C/dMxva5LFWn7e/wxaP3Q/UCTXbA83hrUQEKJTWAXzYu8m
/nTeQvZWiKhFBLS16mpj2XR7fVE16RKVgI4a9O7K8E34H+2wxH0WSxuMGNdoU+KW
KjzVsNf8+0oFAGwy1D+VVyfhsN5qt0IXZEIajwMv+G2CC/fibmXMsl69frtHEbGw
4Wu49ka+N4Du1cTlLCuz7g02bRgFqAWChKvqKUZ9B4CfX6JyPDgUohFtu8PV+b5N
n195drsuk8ZKWOKXO94fXsuq/bXZE1ezZ/F5BXL1wLGpePDQdN8MTqoC6k8zIZR3
aFj60YqfCf1GshIDQhTXERHDC8P9oY2lrjOAjpRxZiBHqW1MUqSFjdVUSEzHFjUz
l6PGN0LVun8wqXm6JN4rbao8NProA1ah2SlzqNQmuJm2sOTMSqW0JEmvYq5wGFEB
+Ht3XMV5z+Z98IQx+Q8Np88eGBAdytLmhkay6CPhWkVclaBichA/+J6vkIAn2q1n
Pf2dSjfhBIFUWsh9i82gLq19qML2mg2PDcG/SKAB/kOnhB0/M9ML465PuHmPkJ4e
8uvvltBNAiIDGMJItCyh5sPct3IqYEPvcZyQ+iukKbw8n0aovF8SHkhQck+xRRG5
jV8nld00ZY17kLyit1gUAzona3YQFoulRrnwqCDZAKO2vMlncdJZbl4jJsvktOUq
SV6Uhzckz4ip/GiThYw3a+u3c/jqivyTOTOwQTzBOT8y1nHY7cGjBPkx1YW6DDHq
M2Mo7V0TURgAcDek4dlXV05l69q1Mi85+hwQBcQWhawFStJPaGSSfYSRFlH0pCI6
4g0bArYGOAS56phLsHBKyuywHbDHe8BbXP8bfL+Zu/98wBZWH9FioYmWoMCAPCf4
LOV/Fr8ZY+48J+ZfaMlYoYH2LXBLdrHKk9R2Ejpl1Tf7v+Zr+VE55aDwWZs+jRRc
EUx4N4EueTPH3dIrP7pakjG9dilnRF31RZrq7Ppvv0eexFJsWTa7BsB8aRvoLW6y
ZY+QlV+NMK3GQOPS/2vljM8/v7StzcF5/a0aFQNBhRI7GScMoclocll24QtdXuCG
mkR19uqXP+tSPjXh3C4Y93QdmKI63gO+cK3dFHcQ99r5SKsllBBq8Y0PoWexXEvG
gLAOGuaQSImVdgMkNK0ub6MCKLKWykERRzLYhnNufTMW/yFij2odpW/YtlSTwm6V
jSPWSGXkC064PcosPNYuM9YhKJ6u9f2T79XNdv/mcQ8EJrrjRci528M3R1Xdfklk
1AWq4B0VloFy/61YgJiRxAgvik1/uGjdbhhxqv4gH5iLKFRxCENCMF7tJTpxtpj8
bSG+cjHXQ2Qcs7hvkzIb6FxrUiHmSxJz5aAQMODVd9zTrZtgh26mopFfyMgjvtdF
4t3e0HjiZNHSVe+epVn+JYEV+0EFgct6jVcI5PYdZomssjD2OWasgbwYSbX43OWS
cp+wuruZPUc4HBb++xjmq2gdfDxCn/8EjIgq53W3qaY6e7JgNwQsYiHKlAfbcIcX
jnIEK/Nk/L5CNIUg+ZIj6WknH84IBgEBzzYOOe2x4vmS1WvTWJvYCWuDRALgOOUP
r16DKdO1SwYgVqzOyTKmsRNdkWtRBl60mLVPVBFepYu2DXk33zmPur0xUnpDueVz
At6viFi8ahVjwcVS9xiSdsmrSi7EC0jLDRnGH7yEX0Vz/CIDcodvbLztxZdbcaKL
Zl4XD/fS94hKeOaTwBpWk1Nv/2IjvJ/zj5URPSNuD761ZMTlw5FJABs/BsRahS5Z
1fgQxHNlfvyKHm4uZMnEbGJqBOoqP15sPdPH09y64BAG4gW0Udae9nzxy0gfzSwY
PU4pZhkCyEB4RsTsn7kGPZQqKTbs40nPE6kWh02XWZs1FEDJsW8ocYkz+s2b/ElO
9RHJNNrHI7pbyBiESTin6liGyPTSR70ET1NWhSI4/Xbmp11NUpMXPSx9H+ZX6ys0
Ubz7VCrVskOHl4B1tSE70q8seB3dYDI86d20oh6J4wLXmDzVYUrDGs8ZmLhY6Afj
NW2Yp/2NJEw6j8DyQvGwt22FDYpXzVxo48gMAZ6Y160VLMC9310ldhApjmOAn5Vd
dM5w3g+wzF5O+F8xBpn9lvlnW6PSkcxblAEaJ1H130gA1Z8EDBraeQHpLJigrL/q
3XZFLrR64UCj1lS19vNYMeDq/2YfN5sqJSP5RBCefqVDQE1mZMqdruDiVE0N9EqX
8jR5olbYCGPyytkPzCadVWQK9Xxaz6hsCLSj+wIX7sZ42GHlgLphs6T7NI3S3LIH
nwLdow0ruTOJa2XIYbIt/ARKPJRwDP7nrbriwxjtv2WcZ8e46rlTc8dyqMygbjkz
IEzkZz+3rFt9+bE1/ZgeAUUhAl6/3XxmL56fUOCxPDWLgS6ttQCMZOUZaL+JNmf8
Mblx3UmHyyD3vhSbFSbORdfAoPxMvXmzGGh7mYnxqQxgUq/sHKEzzhl/RKF3+WWQ
B7fK9DmVeDNQQzgpNxOw6Gb4MiLWHpMIJNfrpOiuCXjhG5zIsZBG9MD0gP/W/VXl
0IK5i0a2bYn2ubqb1AItCnMTyDKEe24AVg1EQ8pr5CtNPi/IARBaCceQIr+eyd9E
YX9iniSGeG/LfNkNN7LZ5rwbljl1rZtyWZJPgUl6LCTOExZRF39ibVePFWQbK8Tk
pK8HE1Fc6gtonHnr09sZiTdHEX77kLWpq9l/bV3Kftp6Uc9w8Fu9ehzJUNWcIWcF
ZO3jvIuwiUmJLDTzsoG/JXj5KoRuwEnFsy41Yj2GXYDxMZ9whCHzCEbTw7IzuUeY
V5RZ58XUNji2PJrj8CEL1Q0rMvL1Gwi3qiz/Kxothu4bdbK2Qxumm1GVJentSltg
RiEcp5K5C98rDosjoHs9GNlOX7v4yNIjHaUobd0EJi6i+JvCOpc4JWvj3/A7CsBV
+pU7YIIs8ns7QEWcfMpw3qUWqwuXx2gwtaoECI5R5gtBWO77LDp+pRxOghYw8opT
v4gS7QWoiQvVZn/hC6iPDJ0kF9MbM3FTNyqATjBHKFWpR8qw+GO3wfzNcmG/YrUD
A8T/QHXaNRWWxookG4NqgqmV0cwXtHAhxZMLriXxSGMeShqiaNWHSbsrlihtppfl
DT7Rcw3m7vc2F0JHKVnrOGbNY4UPMJ7s2+aq6nG9ct8yUxudlBB275JQAJukfffk
naBM2u29xMvcIpv4s7UjospPCU5l29w+cQIW+W76GKb0z5RTnG+qRohbffcrfUaB
HRkD52uw4cso5JJzN6lv0Ph8/42hFYLsNWv1+KOsHDzbpsWVgtWXA540ggGHzlbw
7rzzo40zxaWbaMB60cSCnt8QjhHupgKs64uWxpsK+hMhbbvBS/eK6QhuB1aUbqB5
ilLddzoItHZOr6RqNpojio2hkWlE06D7oCYuOs0SWIkffGXT16Oqv3s92Zh3UEKF
4YhQs9ANIJUnkD0wW2I3lTWzSNfLPfDy0h+9we0TSDti9j25OppCizBCE9fKAGdL
fh9r96Rw9MLKId0mu7UvmqJnSMIkdcPIUnZkLgHVwShpBR0m4Cy2MdzquhebWkGi
8NBFLOW/53E5ACJw2uSWT24lKYKBbeY//uCGfxRGl0Z51Kn3vIN9zSB3a0b2MpsO
DwXncg713Vqi1hlLJD4D2kUzJSZCX48cDfEk6nRKGp1sUcrygbnxlsWDqnAebl6z
SnOkWl0gRuSeoFNFCxX5rq2e9sG7T+ZMqNH6Fq/h3MM+rPohSwL7/D2W3puVkgmc
+G8wH5pu9j2DZOh/sOXF8ha6MWASZcYevsD8IH5NH8ADMdKcszUlZ+yBY+3AWnbO
oR7x8EUz5k5BwdGJKGBx8lwAE1xFfQzuqJwSl9WRk6EcEiB5G/bJq1rJ8MpF1r0V
ERTjfZPxZVq8/Uq/YBsYgtt5BV976trYCXbgafPmqY2hTJZCsk+qeGJpdKswbJ8N
kdduphdn4P+zB7d2vbtyOz4/H39cd15MYkMjNS5bHIMUQBF67seXeNDzT80TvtbH
+h0pciKjmmdQ5Kp5JYO8UoZPWnIXX4O0dI+HYtkY8vQw1LLnPLgQ1vhLlvMnv01F
xP0VKgw/eyuQrtAsznvyyftp+hDM/TgJ3ecxa0zU0GS5TpCGDBHLIwxo3stg9tjP
40FwQ6m6qGxe+PLM1puTyLuzUGy5FY8ItMCafNPdXuqOevSJp1uIQzOgfeVI8jxh
sfTBXMcZeEglOBUh5N5H/O6+yOr/RGKZAi75H4E5z0bHP11TBOZhMc3h9Ieb1zWQ
5KhzpKvrfPSj5E/PEG7CrDahdicZxqDUa5vQQhDIAAStMVZ2nKUytWOKm9yabCzS
OBV+PHffUp0E0Oa+3uLHavIddPI2MofA7F/I5ooQXP6IabwmFR5SFaSXxc2P3tX1
7HuLDjLOk9c20nkvgN9WyiL79b5iKmCWOl1MRWcBcN381HZS6w6EDnniygXMKauU
eJAa0Hx6m+xCQgEPpT0AvcECiQMbUlxYv+ZmU2PkKlSTjiUzQxGrw0PiWQkAyxDH
3YMVDDZPELDqSgVlLbB5Y1qFSkwJPqLlD0cVuyyNo91kySpxUR4n9+5MwX80xdJI
/KIn5mBMw6iSKyU+CzJs74fSYnDn6j/P4sstW2TmUpNrHb0y3BOzwpUZlDzklic5
u9ZfxiB/Uaw0qW7/oZtb7IeDD4lZ3enYc6QAEdnqRULvNnar9Cixz712nuHsReyx
pR81wZGZBkzLFvFA5ydpuuUsZr5se+IpD/mr7Nu1wXM/eh9+9eUZ/36Lha3IwREt
N1Q/16Dh9vA2FGnHdET+19I3TXxE4T+ySxiV7CWEr3rJoK0hseRkcIQdxClV8LbP
h7SPFKkd/GAzFyiGur20nAP+e6qHA8wXEdQHV4lsxNCVqJr7d11R7U0K7tr88Bhi
NyBwv9rQVqjC7HnDGrfCBFHgapT/51hkdL9jnP+L+njVYvvKb4eznFLe6CWvDV7j
uRX4CC06oJ+7h35ONRSrLmtGDn7HLXEiaIWGLeOwEPQj+HHn5fRu+iT35fgz04/3
OLPzZRo+1EHtkqriX/xFX9lZGWSV6DXyGhuDLtR2q/PgAWT/Z8QMMcIB+xjklIwL
DUlwGrc0Xg9R9OxFys9Z1Q9EYUBdJsuvZzZgd5tMDgfpS+coACmvEix/geVpaUjh
G5eYJIk1z8exThX6fmXpJT/KhfVUG2MJ7jQtbDqkC9wJPd1BygwRPHq8iQ981c28
zuZ1ZuJC+egvvlA8sK9QwYHyDRZKK6P/0Rh9ogcpHlWWy+PHuI5bhIeoNsEhVT7b
N+r0H64t8OHgXcLePok5PONsW+5gYx+Bv2PR5Sd32bA6MS/pCtN7XHFpipRRXxUA
BIRWvluxpMAsZ3u7EuK3ctMHykPApqanzWTwVyt+KnEYI3kJ/9c9P1aN3iGMc2Vl
JDNX7nxfgq+VnztinPp+reDdTyG3UV25dL4KAZeReFr43qYy71GpRgadqLqsj3r/
D895G2YKdBUlmXlN5hmjHL/MCUis+9G0jAchbJg2GgEUTayzAMmfiK55In0x7d5B
p601xJrhKo/iuc10OkQTOwwCcyq69IGhGR0EnCnc/f1OCTfEi0IoymaElYRuPbaL
4yzlcsuBF75O2ESfbJwYbtiFrJLXwDSj+wCh28VLMnjJyhl5KoSC1x29rHlPSc+1
91GEZ3/bBWOaD2b0GTI9nR0WtjtQvw70t2r9ozvj28b5yQmEWKZoaBAbRXoJexTY
HpPgdQqL4BYKGY/zTiuJkxJIK+yLoL01U6HZg4Ap7miof0M+Iq2MsV9fCbEy/0J3
RWxF2rgNCwjZ/dCQ1cPZ6O31E/4dnHI06Zi1/yfqvCiDE4e04BO9Mzowk4GoosQU
pAa+iLKUpi7PX2OWMIg+8+rP9onF5qW0oMIjc6OIwyFHxL2ezj/d+CjMh4P9yRBU
g0TS4xTEIxy07zNyT9kFadxxaAC9mbEI8DHHogg2L1xxjtIrAG4pam7e2oDHYOg8
n0nwfSKlAHJ0M2lquCvPvfuqnHsY/TqFPk+/P1pL1gd42My1HrZWwhBZoFSuFB3N
iYmDW2q0aKxIfhAzzjHoUm/pXmgSY8kaeUFbOubnPNNnBY53+26GkQyeamqtHHKH
hYTktxf7ILR+yCwpXnZGRrAbF4JKuCRq8Sy419/MmHmBVpMLUAVp3axw8Ag93PY7
h62fSAMei9PXpurx+uGcD7vGUuBmeblUJOs/Tb2UnEJwajc1PRlu9u3VoRo9rAYR
ZVd8Wi0ZAVBmb5XLdTLx1Y9AYkyug/fu44UGx30+vOvBmVJs/zaeWC3CRWqdexSg
QB4MQYDSlPR8qdnXOQVGQ4lqS44h+TXo+b8UMmtZvmNMqQ/gDyJ03XJ/iHl11VJy
08t/80cJL0+H89d1XbpfPTJM7OQkOD8U+2uiSpyntaBB7SgmtGJgb4Qxq9nd6zix
1gcE03C4fsw6AP8ALxTYq8ddio7nANlOzGzSFzBbCo4WUG9w1yxErBlKwBRQTWrC
wiG//k6U84jHlzTjE+GPyQL4yMIQxZ/vLxwzmbhdPYTJOCoD24DKO13MDRMlM/+o
SLDujaCrF5+grNJRSbfEBfQyjsj66x+8g0R5XVKl0rr/6STUer8jWU1Ez15Cj390
9OvTnktsnPgrP2Wxj8TJ4erjOuYXazJEGr7Dvnl5GYsn3jxLpvDAz+ve7wi3Nwek
GBJFXpbv3bysPvQY9xACNWE5EqsGFjaImavs7LDaXZAu5Di/mRuz+TwIKVRjbopG
rR/2SbxKehF06ckMJv10PHWjrd7FcU52TQ/JQP/V1e3G5rclqOuFhrP0wjfj7dD2
LmQZ4eJ34d79JpjXCH2cEMkrFeYykTa7r4RkJ7S9mW0U/8YB/G/fNSpP+InhVGLB
ss5GZojXEfc7kz/+7NBlRHGZ/jiam1/yjO+sSMX33wjboNNdguiRBsxa2Qp7l5KO
IlLl/8lM6cP5oeWd2x2SsbRJ1r/kJKhb0ErXMSYCzcE9GVe0SR86nyjZ3LQxJKuG
H645Op8PWt86cupbsDUWizgUsfLKxbZgG8wQGf7JNBx9CcvVnG9f09XOOoroLIpk
z0u6MLQnAG2GBvL55cFNTYXuOEafx7FHQbenc7p4i2yK9u4jHUyCxGLf9+qr76KI
myvPAdH6X/Oc98MwJ0SKTXEolztoUmk188NtkX8UMNg0IrrQn56+rmW8AAgncHIi
3iBVWr2GXg/v5DBJbPV8eqzmrShUP0RP7W/QdiOEV0lvd3/WASZghdHVKL7B1kBO
zK/iMFg5W0tq7XLgV8rGqp+prVtJj0WuwjwgSFVe41xWji+o5pMEOlEn/4dBGEiu
R8vBPmk728l2v2zTtRTMf4Gb/OoXJSecYPb9r6dn0WrTnvrdjRwGSFDecaOE+mcB
cbVZgitxj9MiG3dHS+IELCfttHGqOqltPMesSBK3SPDQk6IjJZWLVjaC42u/Hshy
YWfeYKUiQtCIj5dMXhpVa0CRWH8/QHL1mKdLmsgg3lew6BGgREhzhAPNL2QwYKaf
L3aVp4VKBhQU4WTEivouWlP6VL+beBnbYYUj5shHeQawSIZUA7HuJ4AkxK6a3rzb
SsWzlRXqy76Fea2ECjrQL1ZQx+9v6naWEyF2vXYBDdGkAiAd2YDSX1kYnPNQebyA
QnMHHECev0YgZ6pbizUh9mZd6WFQuEokPfuk1xT283C99GWvpmDsc4gqPyoQUW9x
XKUT7u9Cdamxu55OPIDUocqHUkd4kSeNLqrYdJPcI8kkAyt5Eo3vfSQXoCsrgjCK
eFz5jOKOoptB9hi3jnaXR4WkxnU3LHmscvATsezqLt9T3spfzZd+PnrulHKnZHN5
x1k+LAXRJxgO/pg4vKS2m+BTNbBU4CuudJWeBsrkW/zrnW0rhawOHhvRvx9KD+Ih
4OcmOBUBBWjQ/WtfAfDfKUVc2cJ4XtlOFNhFIifKpdx21zPPAXX+8j0LqOVyLRHP
juoB+X5nep5tUU8NjHl/wuRE8AYPDXkSmcZHrZ6S0FHZOvblUirQzx/xxukBGuuR
y6EOYy/PVmjHVKxKX7uHkPrbCT9Iy5KVpECDhtYIR1ooOTxhmZ7oW9dIvWiogW0A
rKeOyO8SUEdcpme+ORZHXlG8p0n6tIJvz/N59sh8OJXbcEhRdW511ZFrhpY/VI2r
5LezDEgEAgkkgSb2dL8BEMD3kPjOy8O8ajBW1Nj9AiFgTQ7VUlG3mpuVIg2nI+Bs
3sw6YyO2xUIXg2qZXfxEz5fIwj0HfhLat7/WjKpIHFTt6+MVxoFtlpz3OfFc+eDu
7pk6eep7kHxm9gD6hK2KKTm5A4jIsP8eTw0NiihEsqZtpldlxOxs2NpXOJXx08K6
P46kgsumxjCsVBEqWUpn8LrDVzNnh5EQ5v8uBmni2JkmtRCmfyILYu3Fjl9gtiTM
yH8G1Cs4ye1R9yEIZhPEjqkV0bvoTLmI4jLx9ZqIQIdxYAQjug26hS1TnIUo5Uyp
aMpLj/Ima1Y2CCUgtkHGZW3lJ2UIY9HOnoPoEMpPxsxTGGLl+X3u/q8NzRzgp/FV
DT3SROggr2GS+BwCNHqaJNJdTr/NtQ1sSFPm1hJr9WxjbroYLGE071Fyd2LxPIRg
dgxg4mMQ9yBJwQbNmXHR7+EhAe43emRgtaAoQ9g3qakjVuvnT9rCiYxEgHPMcQxG
7NA82WuKm45Lm70et2QH4J63gjIe0ZRG5Utwv8B+s3DA38cFq6MBtnWImmFD6H8z
uvB8XznH5CR3/BjCrxfZQVibEep2e0KapU5MjvZBusaChVd746xh3/T8cl6v+S0Y
o6bHtI5XpCuZv1bHflm8BCfZc39yZrSTug3Ny+VwfjTSTm0rrDByHAawsfyHuQn5
nOs4QJyT75IYYKII0jgHk2JKJ7oqS7ELmVQsMf9eU/XlJtiQGqwE7y2IW18v0foR
F0xgDXYDwVFqoL9owIsuVkbbGMDS7AmtbywpXpfsihviCV0xPNm7lPCyH1tfgbMs
zNIXDfseX8u4gM14ARQ4TkE0tGlNSPDqMhbO77LkZ+PS5dKFlQhQyY5Hy6eLhe2/
ELTXsj/N/z150URKTR6qcn1MTwLim/Ktxd+AXBNASVHqoB4Qj+sYtS/uAuGF+bpb
UYONOMBsW0WYZQWjDz0EoK/52+dmByKKHfmtjBURoKz0rHerhjlMrhNX4ZW97qWH
e9N6FsHrY0H1vUGIIEmix4Tm36zyfgNS9Ht8wGeeKymVfOXrS9/SthCT5PdmCZK8
sg22QCCLe+FPuRWw8p8VYT3eC6L4bD8GEglC4IMxOs5B/XDDZIryEweam1qdz5KV
4Xn7vHmDJw6M49w+dz5GYBkK6OgWfFXfRSZnLpT+dmylJjCA8dVMGkdakAPpFh9z
Qvk7z9YUuvdSM/hhSG2v5U3RTO9xV1VLfP2gyXJcLnFsJUy5GAyfVjVZ0kUkYW43
qwec3OOdeYvNfj3iC/KrPJXPZLybNTL3Z2dS21SyyFkzu4l2ItYww+95FZhwa0N6
uC13PGYDYJ7S+XYkGbrD4u5itjgVuWIzhTpQ0v1cN4ICSdgQRY2Zuns9VwiI4GdM
MpgDywROJK6xxFsFy2pd4BQKdLOzM9BigYO6lzrMNcR6JPH1bYapwtzS8TFBaAtp
HbxZjxettcndX3YjWKFt8iSyERfNuOsJuIN1WVEboSsXc+9O4nAbOY+KmNbLOtnt
pcGj8Xr0JGvL8KUjNGAvqIjIlndL2t07tRabp4jfYnve8clCOGaxtp8jHU8GsfbL
DfM5R5qnUssc4JIqWX3OC05j63nXs2EhUraerKdtyD6Tq3kc+dRYFZTSDRvos1U2
z6D40/5FQxW3/zmOUCfBDz7MkzCqU+zHN5POCBKA2rULcAcda6eSwTkCSUeKp9nZ
IrXj3l/HUprBbS4cQOddrdADN5HfDJhVM4+EY9UpCEJSocar2g6aP+02PaDFJ1YU
sE25vcivf/aJNZDmLuGY2t+1N6OhtBU1nTmn7KLRQi7V3iDJJ6hxRGmw8nKAbG37
F57ZCiRnsMF7r6Ob2xpbPhaOZ/AS9RU2nV9CQBDrnWQHnbfqSat3rxixLLJP3Sl4
oAEiwyNzCsMt4R+0vaEk1D3qL+3FZLTnOnaVZ9RlyrqobPkeO2D+aFmMNjmHgunw
41nFq6JqAjZfgJii8aQhncyqDbzeBzs7yPvtNZFrPtbLhL5ECQ3PZc8TSv/J1LQb
wZiEtl7FzyBGgmQHbD+OFe+iNKF1jmvEeJeomQYN3cI7dGG4Cf5zNSzkqUenQ4Y9
Htgq+GsIeWALgIimMWwrJ10vFoRxSVR/UJvlo+nuQHO6QzcdTWupfoY3jjmBoJKW
b90lMzge01LhTRSPwL+3mzbAZQDKj2M5xJmMmMTo5xTU9bQKiz+83juSm3g14zjL
x3RZBxVSSxwCuxljTBtz8qYhYItEhQRsMjXjxNHzRHwOdtKQdTVRCzd5i6S6or9k
fxEpOt0UJA/5TfM0CTqmk/S2LqNeX4xkguhg9dyFqtYszbJHkRvlXYsII0Eqh/4q
Rvak6K5DoLuxiELSrNxQyDI9Koc3SbjXVqzCWXZ99H6OXlkIx4jth/cR3hFke8Vi
cxORkjgXsPMiq+58FTQfd74QUCoB6C+2TXbp4cEo3Xei++fVQp18BD7pf947Fmud
goiW4XyjrfcIp9kShpyHcG9f8f7AtLp7tcRdLhrYZKQ81iENywGJbtSrztI+oA13
S2+Vh9Isv5paJTRv7CFuRsDgZkL3dgRC9jBR+U/AiXt4PcPmBv5fqAof0zos6QOE
g5k2p/r6V5GAP/Wvl06xRg1DPzQsAhjb2OS093j+rov/P9Lmbf8TF9wEBO6S48tZ
lqbUk1ibqgFRfSm4eve3Kia2KZPoNmOLk58hX52m2znME7+nxbv8tY3dD1L6oxnV
jaOhXN6M0WdBvbKPADlc0EoeBzL6oWtWfoLT1l5y2ix2TadkdEKjBUY4k17WMlhk
5U910twVM//PiLqIiSNVp6aE9iIu6CrNNC6cQz46kHXxdNdzCA4AiF+h9YHAV8f9
uJ0he02OLfA9E3iERmXVbt59W9xZiBp968FgpMr6rvT16LGcyy/X2QlufJuVpan3
f2IOMzo9S9dVcP496eV/teLmwJKeCOtv00bgMNULaOypl3werwOQIqvazuTT69xB
OArNH7XY3f0FhS8BpwXFWcM0+FA8IzbaKeq2yPgYZ/8ldVJNypXywIOYN+xe3fyb
yYeuyTJ9vanIQj4z4rD9b7IexijoCR+SxwprLLjzRFkAaoTAyrl+1GL39AXF8Tzx
atw3NEMYf46JE/1iA/yn9Q9EMiix9FK47mce3iJR69cxFwTTkpeztGOr7ldiDjp5
Y67FS02LVadRxmiohFe3tiHlG8i0TyUFogtiPnSF5IijNIAH+7n3i2CQssqxAB9z
O7JlWHjgXmLJB3WLOkZWwsQiOwOFkdMVOx9WNfVTBuzQz+uShQQfReJ6aIHXQL2x
Ux4weoNzQzc6T7mIYHs9cBZPnmXJtHn0Zoso1VaxqexZu4VPigWiEWXM0dTF7aFn
B59tJZ1Mf/eOGx86zKPV15zJXHU1LV70Uo5PyIq5N5NJd01Je339/Dk9x8SqTQhm
C00hILoKEW4NS1YCe2hVr3CCtWJf1EYXPskNrQ0AW1tqhRKyOv/qabLjQSQLrNVk
gk8kPhaskKJjiInGwVEwZV01L95TA/Dg+j83SQie8jEyxDGh3vH/WevFQT4QVMDu
XEB63gZWHxL7yLcddCzOw2fTInqj6ERqA+xj1aMZ5Xw7GrFO6Th901SIGJ+LwwyX
rpBxWD4dqNFH48jCnnU3iv9QgJAsbN3ykH375w/7H7+xlqhYWhIDMaZG3C8hOZ17
FI8x1yNlLniwReSoQmWjcV0awVDPnCeeJAj1SmfiSqLqE8hh/UnAgbtsx6BuSrDw
Aa2VQusZ/sox+v3mB04i96Ahw2rGGUExgpud2nUSG6JPfYk1kZ2Qjy0SsMzbajAz
sINnACrQICrnofcYuvtoiPr4o1p9Pq+oh5pi5khN/gHtgxAUNKJfYH+TYA1yy/XI
+/3GNgHYpxHAb+WD5Glr9idl9gzk4Cufhi59zdHlfylDDn118d93fPZ6+iG2yk2O
FuITStUK+uUc81XP1VMV6dWWWw0VuwC1a7eywuNeMTzVn9Ndn9YxuqsfATMlD/yB
7cn90MQwqZi3u5iLiHiFh0z3uFMkHOj8nLI8YDOUwYpAeVBGMokxFMsQ9hG9s6e3
Fy69BPckQK/aQgihzcMRWhJIAtLXRzkWqcUtXoarXN+XeuNoLnJ508inJ4ZbqX8l
XjxF4RtuTy/pkMSN2hwbuqEmIGK/srWMXHfwDtDd2GPyDme33KdUPZ1N1HS+rZFF
APWgO5s/vG8DwQHmBeeW4f6dhlKtPR9gWymyIc5i24Rj8YSTeFhBNRIPhDM6pPPZ
3mDBqiehXNg0AwVYLdPPuj/prmlprQ9BihPPXaDFM+AwGRmh6rnsbkZSfaCTyBaj
SnCbwQIBXBs/LIgS+EhvDH2gPgb0ZtOls2gMcYVZPVvIfekE9usINsVfON0ibVzJ
pdPnH+Dl5uLrRmmZ4t9ATTvykBxW577ibIaKd3xU53yon25Z+eMOA3zhv66oQ7nj
JB1XJT/YNhwPxCFTk+Z9uzrZSqN2zg+96HFm/vtljh4Xt5GcUEgr2+O6ZTOmdl9r
zSejANkGdp67QrtJ2qakSrwLH3meTjq7fiHTQb1U3te9rkDzNad9eykkAfCAkyAK
YfFI4SR3HL8iYdA5XmF5oCCKi+vOq9c8gaLP2lWcAMMKUqf3+o1WTS9uhbO77S3q
iGbI6tkjwhkJ6qWdXdHynSThLqJerrmug9OshAaUyqCP3UGTyBV2hcIlO2jT1tqw
J+u/8BMfnLKNMP1h7NGoCyvWqpQfsuOAt3zWhv5T7yNzrsIiJTONu6Da9Axf3Vv2
PMK/lZWrdu+/DRcsjr+la9nqDmLBEVh/Gx3vK69AI5vdapS1q1Xcv9bY8y3Mbhup
zTq9ZEaYt8gP1dCDt8WXEGZTbjuYgCu8YqPy0LihhQX24DkCm+TMMf82Rv78KBva
Lwus0A2dhUdIgS1qLqPOfAMuUYgl8FeA3sIxsbAy7DuKxGjWYAZHLpRcYR2GWMNi
umldbm9uFCCseXBC7BdsZ3n6KBPI0or33TJMEgHA4hHovOSZhOkxOetX2R1rT5ML
pAA3v8CEJFPgFXV8fWFMaMQSMnTSXKQvOhrImnlWjjtw+7C9jUJI+zcz/N9Dc9PA
gmbFT8oYKopw7LsbW1vdNfTXkw2acEvH2r5k2Jy8fnCYxHCA+72QYNl94d8eimWq
/BAxHhLVrzPsHzTRlrXx7tATwP73cXbVlYFIlik6CMq2nqOaC6fsqzmL5ghUElLn
Qmv8IB5P4aScW3MvtToHzk3DYocwvzhMhUFfZEnoZyHoXsfeeXo9EHmC+9klaNld
Zsdb37Zx3mZ8oBWnOK5mMhZHtwV9F72WxLBuDaY/6TFQeF528J4iAKa+V6SoGqff
zu4R8OXP5TagtNXTG1m8zOtu4bFhWtL4eYoT6RlqvXJSSjuKpbdIKkZRn5z3ln/6
U/Z6CgO1drXguqV4A3ZEM8qdbP/LIshKwEWTfZw9hRQDAqwv5lMWxKNfKvPZN77P
2AmtH3arzw4con5X98TMrm6wqq85pSxckR+ddvJvmn4EfdQFlmYAeCXoypZliqqU
Tz+E7qnBsUaoSkp5LJ4v8bmfBhMHK7r6QbIc5JfLPGPe9aWaRUtvfzA/TPiVxOiI
NAfu9mRVDL9YPNi3CBEHVOt1W/alNV3cxnLeVrx9wbb8dBvGl4V4amPndE5wGXhc
Lzqr3IzcBjyBwu0V6lR1DxiOLfRMxMsUZUf0ZzeIv7fPu994bVlmr0IV/VERgMrV
GcS9CyRN9wZyIAXIVKo6UcIBJFUcnDYwkI4DhxRCHgsnEXLWj8esCQmGnTM6UBKd
onfswwFplUijKLcM9bK4kA7iRYhU+ROnJ26mmt2EdMpVdjKzmVsbxd26y3dTnrAb
GPJJGYzfRDrIINZR2RRhQ4BpvVK4Nvyw78GGnfGUkz4J6QCZ9qKt+uOuEZjQRAME
RuoisnnpeeExeda/3xkwy6zSDZpe5RfqvxjMkFDmM3B0cjoODZ/U8xSwv9Sq9SZS
Rulu/wWtD2wW06R9P80AB7L41BWPOTBEpW71I+8yIyimKoDJOovKkn8Dq9/WEZgv
FVSCIT0cyWM/kECj8UFv/WKlsrWc71g3+VuUoU7QuEVD1axAMel6ju+q/1A6iPpG
fZ1APdgNWrbvaI2rW9KUJZoYcaoFooGpROtukvuLOeAKy7clAjF6PvRYdd7WBDhJ
pdsLk/P907jKwhyW8SueEvGLg0CLmiBbEejU4LV45cgWbwkjrTrMKYZ3YfdBjEP2
EjPohCPe8TRWdDcXP3vEsAjn3nvkvU/8xL1ADlSmpVbaROUgDomKXgTUrhlEMf8f
mmNK0D9WzDVByslPDm3Kl8ci4YcSek6EUG1gKfFz6A0MZM62wOfPUvAuM3M2tfV0
+XY/tzcX/8kZ4bT3mGmxWu2Da/aNET79GP50yKptB8g4mKxLCA+HzZADhxnWjisI
GxSxSnEU2JMdzhODyQrr79j5+kZdT3v8grnqgMx/MUojTEW4h1j9Ob9DYSTPYCC/
rz2nX+0z5MXkmPZdKwDDFGYpQHLvfraxJOIO9Lem6eQU5sAHTQjKh31XF3supABP
MaTLhHLJ+38Yu4L1wZe9UNxl98xfWtfu7zwskRx5lY5RFOQ5ADIVRcLfn8jttP8P
us9BfYsdOpHnCHjo0+BdFOS+nomE5yhIpFifZMyyqxTCAW0s7nXPhmx1PBiyqixB
2+jCeg1g8qW1RT+B1LvroayFSoJt/zcqVvMUTQl3HYFrC+3I6ZwEgJro/XCX7UM2
j6tLBvRp3HbNm4wK+VNwzWyrDUOOjJIEuL57OZ1f6axMKz9IQRUAGtrCVAZia7G5
u58EEToRM09ppq2UFaqFhIXSWn1aj8Oylppp6Dtem6UbzqY9gXnf6PTMr6Fpfmqj
N4yv0wkNUIEvQvemdj58YbXeszlTBOJrpd0Vv6Rn1HJikr9vUk93KFSxegy2HBHX
CoaXFoGV7uzy531RKjDCsNLikESiYpcaoWwKt/ypIBXbV2WcTGfvwmpPlzutrrn3
JBsY+eut/hMzDboqtj3i0Cg5K1ZhXtXf8MuQ9gj66c24qwST5FnD2BPeoeHKIi66
mJc3l8CASW9EKyBIeQ1hMXtjkBJERjwaWDPU3yb2VmGg9GkM9bJJ4ZDA6tT7EY96
v2E05vd7VyntY3m/MkXltulsrj5IG72vz7pcRI4bbmbNFAELY5sQMHY7DIiRa0Bq
15HPWSDy7Rp70AtWTKFBLnkEyxt0cbymwadxK41H+eqIvfvq63bqplCcNIxEJCOV
lL8OHn/+s6e0fj5i48YC0TRqTUAzM/IIA02IvmI+3Pjs0VqasZe3q73cJMJfm18h
Wdp6w0qaOgnlzDeMIxs4IwAuQSgcjUZdPI0CKQRClnYG8deGTEhbNUKvzwXcefen
mXqB5KqqGVoaMuAD3ulnM+gqSFSnd3X0YH+v6m+XzGf1D6KnOrZm/82MAVCJ/Cz5
xDdYPXNpcRSmScPdqilWgzoxhVmsw7xwPQU44rMzwij00JgAtXvKCw8oi94ByQiF
DsJrr0nY8Bbxj7/nQkWgYqdLQaYwzmpSPAhSF7FJRsvfbrctE11P6Zwl+ucbjhSE
RLHoPKdsSvns3oqgp/OjOVTEbQbMzE2BS1G1VADn9yptqO9BhI/8MlWbwojs1hFT
InBQ6OW9R43xDxz37okCOMELxxZLPJwP6Zyaz64MTkKi509514PRNs8OCVkTfrTx
1iYFvavsPJgGcfXY2TaElN8r90RJF68Y50N2i/La+Vc9ag3c593jqYTi5/HVkBWI
yUK0WIET+TTSWOdmMg9bDgZMSnNIidWz5CadftQFMMo0gXLNNy2TSwBXSyo/IyH2
usHGSzdZbPudhNZBRkoDzCARJ6OT7DwqY3tuIWIYRgO+euF9fZCX+YP+Gd0V2ohD
tuqHLIn4N1vCwEiPnb/1hH2As5cR38/F0ZM6Q89nJiBIvpOa4ZNtlcdgAawE32NA
9m6Qi/5Hrw3XhejK25zkaFVtrJQk8lgLaKie7u+LqjUmq/kq5zGtoSpuHj9ri1mq
QeambTmDUZE+7ICBKMh1bxdM8BuNvDdxXBw2bAS80/R/tfoz9pvq0Vr2VLAimCud
jkBOEZeBLd1jZ+eBnLFjNA9ZlC1WW8xXT/fde5RoQ5wRVQVHv8UezkI4pFcj3h1r
5FJnpfuR4Pt408d4GaJKgcHDcowkTrDiSyA+WD3zQPCe2AIE26Mf2Pju0ATmsd5Z
Usnz/mePhHJDyQnldnVcNJaeu2rxWn0txdfn5qofkn1IGZ9Ut5uaEC+Qip5iKcMu
5wleQ6tKMyHTKu9/b3XW+jDIFJGemynq4AsGrLiSNk6kcG6VrHSlGhxaAz2LNSFa
xbSIazyfRT0rwjg79MHlBWTM7dcuj9vbgZolEcY2MfgzX+xzh2+fZoTnIybD/xRA
1PiWO4TB2A2T6ogohgWcQrNs+VzKHWX0BfJp2cYsWVpTL4zAyLpQ/DtTTGkUXBuY
GSc9OITu2ajNj8uOgMBDLJz8Fn6P/K/zqsBOJTwkGHvtN6S5E/d5XgUcsX1ozlUc
xbUgrwQEdpeCzhFSWTspEKGkwnUqcYOtQTpGSlMwolDzB6QOMFYqQHAPbce9x8ja
+ZTQcqqnvOHwpF/jsO/7j2GGRHgjeaMV4x/SyBK/ffQ2jUD5JWS2LHGWfpMEe9lr
oBF0tzXeymTNKDOYfTNlB4hn4ozD5eUDyiYAT4GXaaUaNeyGFZwsU7sbs63ZZAfl
2I7DZpFu/sQHooGjCnf0G3g75XNNb/Vce7yO+U/CdTfDVCgthPBV1FQRx0n0aY6Q
X1N2Ow04fWQQ7ofVh3B883mUg9Rf1kh3LDRuxA/Sxs5wjhvxGw2yxZMiT2ha51/c
Si3mnERJhEHQ+AetCBfnlQ2hhwcpYeMs3DFHFFhXsSLk92JWVayTCs3Pwt/7VKw1
73dfYtWv4JvezqWxSGvLvJVf8hUjR7jmcJkJzKHITUfWyz1Aqc+zw8ouNEvIHY6A
lMZ/37a5o/1HQts80wXZLvqUGg+UOYtaHoo9tZ6tUoXrQff4b8SDqXZM9AZVn5Zj
70oB+pZRGXcXi70EmeOyuE161TkhXvbnF+WI7M3qcKNIyTzvpCcIwrfUoCBBC9Ld
kQMfvUNiE5J8tB7a+76baDj6RKAkldnE3wE+jkPGkW6snbtjlqXcy+3D/SBZ0AHd
f+7WIDR0i0PhH34KhfzfywHaS6f+gbfoY6Ko9PExKZay56ij+kxLWw68mW3uYLYE
wXgYEd/sSVZcBrE2k/qJYYnzR+BE9rDHAspXcXqILUuKxH9NBfH1SlviqItIBZgC
SDX35ax/EwyhyXtMcNG8ocYYbZ4JisvS8Vb3+KsF/XRdF9r/ZZNeBYWAVMxbCExD
1dUkWmNgml7RcSNcaQxI/Z+5RU0JThP0o3SeQxxv58EMKM/dn1pnjzi05demLxN9
1zSa/fq0VkVsSAaoLCWiGOgIcLrZqc+nA00znH+zLmgqbPiGTP2Zvq2pt9wf6Zox
nhaoiwgDEI6A4uSd47TPMf7jROuiGnxy8eNrC6SxNmUC3U57xzPCG80jELJrqYGG
+HTB5wi9Zd6IGNajkQML+ZqtuMbuUQuGyVRGJhk99aDsUWl7sm3oH97QsvgVc3o1
GNOLmEV4JktMu/Ozx6JNKm5hXttcUuo7PX0NZ/V5SWlKjsiDUIfoyIhKeThZJbbn
gmLf69hnyuWNwLHYim2gtv1eTEHvrKFY7DYH8yTy/qpBLELCXwS1c3HLr3ehi3zw
kxEcJYiecSX7CxHLucR08eLzbPbaQSbT6hWafO/39BQ/xmmYh25N+FZ9inJb1Pc0
rvGYME0fG6fAsvwCqZAMMLrBvmSKUMH/x5LKdzZQuAptQ992s7jhPm0Ngp9zP78w
sjK9kqifY2AWGo9bIdtg/mYE9kWYZDa6H2yvMOnvifztwf3ipC3XbJpefS2O0olf
VlDQX9CY82+N9NpRvbfELbQmD2XVoSXZ8B/YZqZT8WeFjkKVHDdwofWVSMkgCFvx
OI1BQYJu1gJQkrac6oBsobTuACQcDhMFko89WznFCi7ZLANsxng0lnGDoJvxYf4/
zGcqqhDYkZ+ZGbNhM+IgGbFNn+pJcYnIpbnWYPJqF0nVrRsabipsFfJDkOa/09QW
7ksFt6jQktBhtPeLLBIQg1hiAoHFplAGSKyx5EkLdCEE5m20dUoNC0Iyuj27476h
hGTrHrobtfEJXNsho2a6ZQ1IukX8TS7t0PVj1RzcZuyxAjrlkFSWhnUlHdMykjbQ
mDzYTpRznqGLXBOmmJ2gSk2MqTZ25Su4UKRtV9Fno+z/movjEhWi7Yck9eC4VIw3
lVHpb40ODWD4cWmJr3DvVIUuZKTOaosj06jJVRzxo68gtYs88wEzcp5aaSinWu5G
jXb5KMcr0hEZV7s/DXCtuAryqdvV+QVMJ/6fEU3yvAKt+xzbTBmDfHyM6+t5zgow
3pM5nLsKPkz5GRsRLWKVAg9kU/yyBOHsWKkJGSPv8p1meNfYGjosNUNQruJbat7k
OY7q2Yt29oW6URcNqytgFeXcTarIJ/y+JqWPBi5A/+3Hn+MNxhJ33DC1kQ+WzppP
TSQu03fBjeU81CNLZP2l3O3bM1BWlT7JcX2qcWr1g2kkTOvDBP++R6kxZvWnHnEX
MWel8v75rWnEUA8c7dZxWxy51N+4pRPHIrhghuB+L5xsIuBLKgoW81Td/fr7fnyu
mWR/WgRhPFN1mFWAzdexk6Heaj2MzRgwKV5LepbuOFyq5+fqFP6F+bRQgn+pJD/+
fQMl8G7ts7V5bWTTruLKsAbWmiAvwnBjLQx2qNkIcoOXfpjDWWnBH2AvEdd3hB89
0JNQLtq8wZpNfU4enZilq83U6dY2twvpFm0s+Y+tktoVToDDBdWdgri0PIljq5Gh
rhuYwq8Lir9ClgP3cTQrT1s5YyD4cZqH+CQRDghakQaYpsvBKEIGph5ccAPPTEjj
qj+0vEfHrIMpDqW5k4NjeX+1azVFt+W70m0daNqi81TzljesaeZCANGGNCCsKPEr
U0ocw60QKBoMs9hlSKVAvlOJAugex/vUnSTuOG3WvDFnu14cVMjT4dBATvbHzm9a
LLDPyC86M6Pm1XHxDANTgcHsdZICJpX5vBPsD2ioxVOtOVC+zXkGPZg7rwi8+W2C
ZgWXXdLBqH8M3Lj2Csz6P6i47KWt24+H4D4F8K6e8+J/IFU20KSXhzyLI+vEuQcg
TgUwmvPukVcJqK2NgSdVNKpb16MIWhkhaTWI8TB6JDH6ry8n+boudapIY38p890b
B890uZOptCdJ9O7Ap5n6Du5bn5FcbjHUAd+/6T/DzBnMXQ2K3Vl8nVLTX50LfPGQ
2dTrdplI46U8XUatSi7QrujTXJRk0Ho80zAwjE7/NW74cX96JJC/xnAAWjRw7orX
SH059gTRyouf2UdNEryws3mGFvTmD9BThKmz8GJ5hPmbKXktYTeZuoZ+JHohWEsB
1nJsyzRf6y79oeR/wB3/0eqtlCRh3mLbhHaxMdtd5OYyqp3foymuyO4vaWFr8i8n
/6Pg3zB7DO8f8I8CMJdwABy7LNVQq/m6Nq1RFoOl2RPFHYyxq1auyQDUg5TYT7jW
enAlaGu58C5sMgK9UEdqtYTzbDZ5gdfWanvcxm9hE+IyVfpG5WLQ0NLwJuTFELf+
4Y+sO3ROzbB5TKugSasnf4g+JTMMI8s9KCRkBUc3BHjNiaBvma0GDJjSdzjUBdwp
o6ymkvjCeu5kzTUgdiGJ7My3R3M2LWFAYQbxFvvjx8EAd95rvufhenaR423tg23e
o+Whi6UBz6F9WPzDrDHQHr4Mpn6RmUJto6SNbTY3VrA6EGBQMeEl4YPQYha2oEMe
FruqO603jlw1z6LUZ2v2LcmGuaQX2aAeyEj/lk9cEEQirqVdtcPoYt4zu+aQH4TE
85+2Ur6p/gaZ7l4Ibj1cvf5JYhA7ltowTw4aKQk0ZIiKm4kje8Tb45nQ2x33c7Lw
jpMxpivNu8sLKG2G0kJ/njuo4m+EkFbsgLkfVhTJdiSI6NC3EG1ZGzfctle/+HQW
54hI/5GLuxE/ioGAfRPAVBHsHglXUQD9SQTFJ9keCrfwyWGWaqTeczhiN2ko9drn
Y0eB9R2ZekF2g8B8shIreBm0q/Tc/UVuUFF40vDK2GWd695MC5/RdTL3whlIJlH+
Njx+NRiEuGhvpYFt1Un93zmcrwn0Ejaj2VBEYW6Zrm+7IdnZiPA69cSNy/o2LJkq
CJ1Sm3SXZXiziAUvJoc5J+EoLQKoKcqr79WYhMEUCJyXfiApW+dS41BA/Uxix5x/
wn/5ge232DQ6ytVwEOI1TBqTyGXJvBbfex78QACd8rRjLNC+buIYrp2lCeIl47Qf
qh5P5cP0HOZX99rhBKk3iKnFMimvFn2QAPtWOmng5Oep7S0AnHmjRPbLM+I/0sTR
3w0TMSSA1Ju/b8Iitx2W/ocoh5+a1iYa0LGYSGPus0zgF1cFXYA1Xp/Y+6wiF4nz
oxZ3P4Kg0Vnizp3UDqiC9uJcArf9u7nxWj7wy7zF1IuXJckPa63vVwla5ltFY++C
tzXc6Nk0l30xgz99gy2GSYlX9ieSH/CcuSGE91fyoYk5Mf+JZMve9mNCOSI2UWzb
qAHvKsJ1h1esVO58aOsClf+HwRWJr2qhnMNCYlXIsyoydygn+2TkVV9RSLWqYlNl
P3gN2yujOR6D7KWWl51Mu+8U+hvQMZjlCIQKVbYAjjA8DkJgpbCSHYqdZUTNs5R7
nHJ84FA2Bd3AU8+SSar3EV/i4jiq8il8Ckb1dk2BnYvJIExEKOTVEgF7LBIuHLGj
aXBukR0x1B1LW9/Mmj9fjo4KLhDxXqQiF9ZYGN1UTPbOKIPlPYpXaGFpfN5SrDn+
lJoO6GWQEnhXlTFsfPg37y48ZVlkyAGFKMV4CxDvJUBK7eaXGUL437zIv/iCvo4z
aDNy0vifVGYbTVdr/iraTCEkpjBEl2tUAPsE2ExOllwexhLg7Fen/da/dzs1KdgZ
bKC3IqVkhAgbLWS2Cp+i/7CE9bwY1lAo6FUopd499E7XukY4FXOnF6RbFx11c7oS
LJWC2Fe548A2R7qRe9XLgpgKxZQsEdWNtbR9VnmWwZjtQ3V+QEHVxk8x73asbeaz
ZPcJFpWcrOICEhOZ2pcdhoAsPy/v7sikF1pURLtADY40qdPpwIzatP/LkvrEIoRM
MbjTXsWSl+d/5Sx89vPzprJvhQN7Fuhe/KVkycgR90MFiZlHtDyJLmloH7UBjQpN
0rma2HH4/NUsD6SK9eIPoy6oWqbwVhePDzahZmPwO7Ig23W1paBpldaFaKIrVpeE
cEInEA/gv1ZZa9Nri5bebZfKuR5VKYTGTB+YWnU9v7frVUCeKwmM8oMX3XTj+Iz0
m9He8AuqDV2Opo4vCgxOB32kGjz40f0C4sTU9l/f34rec93d4xdaGt3wey1iu1qw
RnrXQHY7s5v+SBEGkg4MGgsf4otY2XnUQwGr9tvxfV5dvVcsrurZH94JhKkWGKJa
kkac5Ndzd6+63rOazi+K1jLkNghqjmwuEuLZfOo+osiqnf524pdqc4FocNjXPY/M
V65kqduGp+lG457GVeMGDnqF5htWTwbDVbUar8eZhwKI7cbeC/Ucrdn35eg+zzDs
mbi/7Oq6USXGG8D2mJp3JTt1HK26Og5oMihfeAxcnV3eJj/AQPCUyfbV29pqh1TU
omS2V1//SLU3/UnRnFcjf/j6w+SSsjG07tMiRsmGWWtxcbOfWzL8L4EEG+p+r0Qy
j4GaK3balUCXD2WQwxHqq3Wb+Rf2qbDL67/xxSAiDCzrUw+RZbsjBekACfPZ+D2o
550vOeg3LZG2JApHw+Wz+VZnBk2rf4LHu7mOGcIcMM96PhGd8tfJybz9JXL9VDtV
Lr84a2rUfZw7HS95jtCLLdvqrgKNKFQAhkkf6R4mvnGs1DpIgFiXunf22spdQgK2
X6EK8Rhg5XwpOJD1JirK+fuUYg+54rNt3amirDgOKjmGmHLR3FJiKhnQv7/hi907
OEjfJ5M+DVx4cCV9sQGtfo+ttvQ59yc2cnJk+2NL882/WxiSLoBtRRgejGQH2QJv
jD8K6IZXn4hE2Z5uy0bo4cK9twdCchSUvkLjL3fGe9h0Kvr33hlWRPA70285Uu9o
Yj1t41yQfVhw0Lgu9cLk/h/dkq4fVpnsKipKp5QX/U03jdDr+ViZsGrG4DUsyzY0
Ulb8HQz1F9dE8t+0Fb56msBrt/U8yT+XTZTJho7+epb79a+55xzIZg5pAvHHwMhn
naLF7hP6xkfSMD7vfwfgeazT0/cFey7F/0L5QVE7vLA=
//pragma protect end_data_block
//pragma protect digest_block
lk9nExOm0LljwWw/NNkD09KUocc=
//pragma protect end_digest_block
//pragma protect end_protected
