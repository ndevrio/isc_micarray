// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
q9Jh4rj9yDyJA4qK8ucWMSC9dsYQo9+Qk7+pyfSqsozmdpYBRtPoKvRAn1CnOIe7
InmKRBNht6U0CH9xF2ssKLBqe4WmM9PDf0XN5svvwjekpibqjCblfNUCD+f2U+8p
OnKe1y+V8MorXVkreY4892jdsWzuRc8X/RfXdX+JmNycu2GoyrMVYw==
//pragma protect end_key_block
//pragma protect digest_block
u4rbnRCFLqI/DTw0Q6o+Ho22Pn4=
//pragma protect end_digest_block
//pragma protect data_block
yoDHBwQFc9S7MYRrmpB0TQwv6pPRizr1jonLCDrYNfMbzu4fya8idzYRBFjwnBfT
zg6ghlYfnToCAGoeaz84zPhqTlt4/QrJ/1pUqpLXXJZDfuKfGdIRnVpF3ezcOdJk
GPGN0oFwrydQnQWuRkUJZpsSqSQDil3vDWZUpk/8UtVxFGgTUVPSU7I1h6lSjQj0
A4ygVBVnZlNIVuVwO+FhnIFjmJwpFBhnnw+bUrRRfv7PluVhl4Fj0GgmpXlM1WvC
mnHyq4GzAcTxjBOMxN8lWQwEhQvtjAHDoEicCL0t2CUi6w6baazaokyoD75DEuZ+
F517wy8QrnDqShQ06S++ztMQypGr5J6sh8VEE4gXOjVlZvuV0Url74zQ/YN4BlTI
1rCqJkOkAtJaGK25E/Bl4NMkUreUTAQ1eqyMJy7t3eXVp6qqAfV3UtBPscGE5fje
mLSiDqo5+zhOaNBKRTZ2lwvteAkOINa+bqjjnPVENF0WMaqMr4xh9bHlHb2aFzQF
llboGzmRVQZA6IhvZIPEsXuJ4g71nkAyhyw/+WL/8dyxFEgvvbFAEOgR44PiJMBj
YPGqLAVdcZ59H3D55nKG75Kzx7uxYzpoJDGUIN9WOzWC9ysvNZcs612GzsjLBwNo
cb4FufFeQff8/ujsmgAXr45m0PDTOBp79an8oJqx5/loHopuCRf8ukT0SI6K4gci
qM9TupbGE6J07J1RnKWu+Uf7PUQI2i1h0Roma5RHkrztuN4gwjzq7mLs+2dv8W+Y
hrWnsE+DH3W3voX0nBCfMVYQZZp17oW1AxpDne8UtgSDumX1NFE0K0AkwGGR/U+I
CmR+Fwh6i297T4zPyvojwz/Gy2RGCme4mRejn12p12U26FbIIUXF3i+uMcv1dbv0
OlhtYJcFWRtKhtO1DRl9PKGLg3e5EBBkaShxxEdsPwgsZrmd9iqo+xqG7HpiVcTD
Ucf0eJE6OpddqbWkoU0a7v+8hGpBlGPZQDmjMlOmbZCl/YhZ3y3eXsvL/kH2HrpE
ENe2tm5AFuquvhDb+zSwbweZOxac64neu8RgmvI9AsPYC3ybtg99xaxghAb4K36Y
yvn/JTUudZXD2xIXVsE3TLVOkV0MsTM1F3E7wcpbfu++Ft1mOzoYQT07aUmDjzF2
Gj3Evb1sc5iA9Rvd5JLzyG0QVZxqQaPRLXMV8lC8wRG6rQAPTGuRpj2fbWmyRcVA
vUdSne6+6whykFpJqMxvCJHGnfU1LeFTQOa3czsGb594eIPNh/X5P+UQ8ljyARtG
50w0pxRWPQCD3E8D5/5GMEXC6OqBijhcap166/I5WcV1o492x083F0+G3oEb2ey+
TPdJw0U6A6K/AXHdDzxcZRPVjYNx6t+Tu/7wY/RnnUVCglRyoNcvrOQxKcfEhhnt
BSZS1jz7E3/+S7X2mG1/8CvSqooqGGkopLhQ80EI7WlttY6F8PsLoOAISOBip17K
vrJPFR2oBEGYDK43WpnhkmMGyXJTGktG9oFlvPEWFpqMQrehEOihnTMJMZ7scWum
fgxdWn20Dpvdyrn0PJxtLMk+UFdTwOfLeKjRFoITtla161kNrm4zq5R7vBi1NTP7
DNOVxdUfm1lm5LC9QIbDuNmOHvriiGjkgTnn90OvUefPXn9gWuMTXBrywgAHEccs
INt9hYl+xFVlaDPUomK7KSAp7buy8RKsCt1SMUD+AdZUDa/REDJ6rSXnAjyNZANl
HzylymaJ/qVFtYEc5J9RTmBDS6544mrEwORH6H3ijasa9TnRM+MSpwU5XbQcDlJz
7700LimtSLucQX44L7EHYTwwDCen4n67kBZeOITewwQO1nvRQUZDPvOLYqK2RgsI
jIvLVvv7YjDRWj1Ab6Q/OS9KsGbosjnAQYtcfKfHxLvsH/dymjobz5VCX7aGPDcQ
uLC54OUeowcc01/6UJ3MYjbFipn00m5KzjkrJvVrDGe8iWz09vBkW3nzEFskYVv0
4kRklf6LJuBl2PmBF7MRR79n2MIzByCsUH0JWQX/yep2PFjon75+BBpIMl91YnDP
FmSbFegowl+PegMQNWqgy1xdZPZK2FdmM11mrgy5kRMRHsoWL2epxrHY4y1lKfWG
5CvzAkhvEXfnuFRBxL0M3jrpxND5/N7sqGhzlvE19RzQ8AqMZCV1ceHRG0IVPJw1
FkfawUl8tv1/3HoV5tnv1ygsCEyxQ/eP5RsdooMl3wXAZ/v/yXGa4VRZrTSCrPlP
PEj6VzRdfAB8wtVKhaYB6fyN8oZVn/UPQ0FBE564ABEJDbLLbptuTdME/A1bX0A5
WXhWeRDcRZs1IA1nlcmuILHLjilYKAP1PFMK5+hCjZiXgGUCccgg93nd6Moraiq5
IDkoC5GqXUBQ92kRbREV5Rqx2E8FUpN1lByZtoBIPOufyZyCeM9wr7MK8qwEsdP/
eVa+WDSIbce95w7r9SkDa/J/tDDTizzStERyASaREwvkOnDcNhGj2HVpV19jSSOP
8L52U290BojQr8Ygz8wzYB9tKHSOvMbru9LVfJ8E4nc2NHeRsfN4Atp/vb40jG1B
5sWnl2ptwlfG5oLzztRINNT/u5G+7xPWegYOnQeSoLawl7QvfCE/I4P8idXwFyh9
7uUV+TxdojgHzieRlOd9Hp4vqFo/IBRWciZ2d+pxcSY9V/evPAlnWI4XDbgcMSqw
BMrkxHOUjAiNTzd4ZPs5JNy3LwHJCpaFky+YpNbxFr6AG/ndqdQ9hI5cX/eBmA6S
kwBXUwQB+mc0ogJO4NXBxhJkFR9w4I7jM6xJrh1Nfbe2UghiXemVC4zoSPq2Neww
JXtPsikqCwoN9+C8YmP9nIDycNDMzHQ6TSLLf8O6DskitIbTSz9KwaMYXwRLR7tl
fB881lykTVqF+lDt30+OzQ==
//pragma protect end_data_block
//pragma protect digest_block
Zra/4rlp/OeBMHhMxY5sA/0ZrIE=
//pragma protect end_digest_block
//pragma protect end_protected
