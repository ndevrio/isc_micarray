// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Sun Sep 22 20:49:28 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
j7tmn4KE4uOZOVTtQVp8Fta9V9vqiGtjmoyErS3XJJE4D0SC/4q1++MhFJ18mm/s
LK0CXwwOAc+ufeBaIKiX27GuwfMcrhWUW3vXhRMNGIaths5bIchgq+OYE6FBEVKO
/zQtD9DP7F3+AekgSHoq8XyJEb5xGG09znV0yKhqWXk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8864)
SNn5k+jtaSeDREOJdYw1x0SXUaxcO17MsjSot2Ft6CaxXdsVEsxyk6sUYxJ/kOX3
nu5uZrM+GCTy1FGlM/ZMgFTcP9TmuhowVAZgFi87Y6YfVmchosBqrDPN09sqSHNp
Qn4gV7HAg1qAp63kKxOxMpj5SJ3fUK2LY+hDderF7meEZKFnkXGZOodnMGNTwl3Y
apeY0094uDPrX7QKFGPrDCteVHLKQ3s1YfMtcxzhov8net5Wu7k+vReqvlYZNR3l
nIV1hxzsd8aAPXPJ4t17YIr7XnWYDWYnLeE8FrUiwV0jcqHlfd+CRX73uvRitpuJ
6asT1XwsVcTW5FCEjQl/9NcxvZelenr0zM8s7vOWPXa46Zf2C8vLsgDyPS+czh0E
hKvLq4lMitro8HAvdWMgEOX3L8YKU+graahUkHE1mAo0WzQJEq9TgaeuUiLY/lIj
G1zzJw9Td3/8+lAqHDWp+MGfr1v7Fhb2iKrTsqVsQbC7Pl8/gJlrVEp5Lku/vjPH
/hayaE6GCseqzg3RoQOVS8rmPjQjfXeH0QHM03U/vXUEp5jpLTxrCUpklhvXY2ZO
pyMTenwC1Vd66soMpx/vYTGry0wulw2hlW0Qw0Q/edf6ulqG2JXCFRNwoehRuaoJ
3raf98SqgBbXzr4dZoRxtzz9Gs9MKaEasOEmvg1A68BnzoEiwfrm7f14egFErNxk
SC/8roQcCKMFHkUQUlLnSjrNnU9i9ouiB/hm2ZH6h3NcJvKEvvx6fYPkYIjRyUhc
2L4Kn+yJWz1oEYMnsjuvZLlnIn4I00zkdVIDQRnAk+pt/lY2VygFKMJ5RONGhxGc
aBGZZZJLBee2qamnPrccXEBcqF1szCabafhoz7UKzfLXLFOtwnqt/KG84uv5RI96
27PX8UiZMkv7nBhgW2FI6kQtd8aAuvmGfDTbgY3YsAgXIciM1P8VUw+cj/bo4trL
7LCW9E6ZszrdP4xfty90gZKr/ZcVa3nCHdl7wL2ENcIqqZQQ6lwzfB5nISOP4v/n
Mmbs2CT6xDLHb+1vgCuHAqZ5BIuKnKyBOCCgRwMlp5A3NQll35MJPE/UIV8KFDt+
UEHE1XoIN/QGWTdPK8/4zoA7M6Bg38WjPf01C9AcS3ngblbRg06fIp85fSaTS1YR
NzIfj+avxQMMm9OizHD6NFEYoOvf9RpV6XkqcK6xPv3qs2rHMG5CW2zxt1tGifAt
4/nrtiaiv8xbSREGzLzrYLWDaI280FInjEHXMPJoj1KzvKRhW/ymxh3ZFNiG8yq9
PhZb/2O5tTTIAwR9BDJ2oxZ7LlRLcKQEClwNVWNbc7tAFdn36WjLKGYGgGUcEoXf
TUKEqRsWRRRCSumErIep3uGG9JCs0uuJKyY52ppeCOsJT8NHAhaKsoi4HrK4wpeZ
jIzb3Q4bvP60sxuDS3ACE/27WmB1zQz03TczbFlC+n6oyUiRCe2ySve4/0q8W+T6
Xqu8g0KfxfdlKWPK4tlMKD+sIbDoG4gI0Koh+iPn5+Ow40lim0UlsQ5vYnn1emez
pfHMH0uD1L3Q67prVxV0neH31dg0FkczJpvh2xVlrfbGSEyDq/OvFtRHdbvyh2Cs
DouKb01Q/s1F7g3PgCGgNOABHiNz4x/iE2P8Yk6Y3utBITVl9v+7UrpTsfZXe6Hc
lN5B6Da1E5L9VfxYpC7zDVn8/SVvHZvvoOYUB7W8C3TjqFTkqiljQByebvk9j11w
8t6ZQdwLxgkdLavUnqi6kk84JvY+kleTNcXU1ypn0dGhuaOkfFqMpI0KD1rM8/vG
43zw8HI9Q4Nx7Ugl1FJtL6K/dXlbqHPl7VVqfXLn3ziVbjHC0iMCWhqXvgSW44dl
NAhNHOmgasbpTvioMKK/HYKUVtcrTYrDr/NpZSy158STXJDo+m1B17fC9i778Lyn
A8g2wxadu5t7n3L5h4Nlljkbi56ddAZeTaZ8l2xCKl3uA/9Ub3plfLyvUhzhmQgQ
hJVmwesV0bacNMzKaD8c+0bG96d1ARWj79Lyt9VeLPVGDQenwF9WU22Rr2I63WO8
37caDTdQRgxXgmAizamrPthxaBL2yzw5vnNzKVuxz+5S9NfHO/CjjTVB9mdftOQT
9qlQNFkCaY/Ex8dqHPbgzED8P+3SO73an8A5fS3KtkZHPnMlgpbQBWYA3J39YBQ+
sG7916Yqpih9aXo+UtaohsPKCz4Wo5Dmqofn2x4EnwY9VGfFPh8WBBUAAdFwi0UV
djw+OWjbXATkfoUUKwAULPNQRTM4Mcim+PVzhYa3RqCTwIgcZfFxZCzqLO+tk1j4
O6YoRuVSYIMIZpIEsaSc8LrejHnyg4QgECR1FUoKu7s4K0JaJ2pq+t9jpJ743W+z
S70rM+kRYOTa89DlP87EJ8cudiN0ysRBfBU2M5y07pR8mIfht3tV0aMfYhNcv5G3
2GnIL60LMbuUjEb7qqjVLqOwTPlgxilgQA83+wY8xes8W3s9ywyJJBsp4Q3GSfZ+
h+BK1gDx5fR2XXdFuF4NvqB9GLc4la0gXAn7Oo1QC6lvvVLJ4xyY/EjFOAf2Eiy0
PwtyBqfHjs1hSfHQU+scNsu1bo9DCQTZULvV7X6291d+FHqchorlXhpZUwtCbCMJ
oxJ1eQ09SR7+n4ogrVip4Xxun0jszII3LVIIKLegxcvTmi2H1OfJnwuoygilMIgv
r/JZ2aT77O3R44A0qN2GEEQ7wxGYFmWtf9AX+6kEtJ8wfKC1m/tQ5mpwVTornip4
80EylIiQfBO5lsaaADq7orJbWO/3BT2tutgswnwVWFJlawT4UBRq6lKR+8TGizc9
+ZbyZ/piyPzHy4YZhetbIH5/1/oZwFGCSI+ir3sBjtkzuh24KzwurTvZ+DnT1SU/
7SUxIWb4DJiZgMP3U7bNWj7JGbnXiWjZlcv9Cd8p8Ikd8Yc/VQGuywt0+itW5mBF
1thLUVOQzcysmq19wAHVB2oJbw41SkVwKTDQYvplqEz2Py5HqrHKXG+nzdIpFkJH
uyyVgp+r73lMN7Pgu0l4qOmNSzAJlLRG6ZGHUQ0LXWVjwulFv+QZyJcdB750vK/4
7y+rDfWGq8cAEncdKNxNHXwMaSv9znHD93ny13YSge3mi7BCs4WQT+NxWz/pKBEW
Qy2B5/Q8CAaOG0rV5FUnLiCGz7qZF8Ef/SOYtBwkFIN7QfDVwWS2Q03La+GfxWEe
ScI3rU80hV0PeSLHyXN3STfWSMqLN2y9kSdUjTVeULoxlwCFk+tf5IJ5jH8O/uVE
tz+PJGqzosQj9NA8fe3G9rVGUVMqKGecnPi8W7DPJzmtq1SzNe6GH+nS4+M4uJre
ySQdTZv7NRpd2DgtNzQaAPldeHpcxysurabPEmqal5M4+lq4kWeWaRAVjYETtfM7
xrK+5b4r1SnHkGg9tfXgonP+HbRYcTEdTILIvxAaPZyV41rnSAZh+gocIMaaMnhQ
K9ngwjpkJnEO2mCiE6n7uDf7mTDjcaAeS9vPFT3prEJPG+5n9NkfCq7NxNw1p0vS
7YIgzbedB0EsW+futG7H0quHAU6h3ozuZcb2SpoPW4ODnsZbaR4bLITSRb6/S4CA
okJ+GITZz+KGQfj4iSi6vt5MYo4uFgqTM/tVwCJK15fL+Oyjwy/UkTTqg4Db8DRU
aO9d08VdYLeqxOenzlSoXU5ckjT2MFRGyCsa5Xwwe7K+Gb2Q52LhaDWbpUjWkO7x
WRK+FA0C4t+rEug6kULOPAPUI8Bj0xQBsfZeBKayUSwshxUqacugM4pK9gNvDjtX
8jeU/IX74zToEeC6TJ3sEyKBUIMM2eK4VPGdR75y4EPlBhojsneyUvgSCIFLIShr
Mv6+4NUFowjhJpVhoB3IeCKmOsVahNg4EAYwTYbkwZiACy8CJ+hhKwTgC4gF2Cdz
sJbpYHyKS4bkMhuAf1DdANVMzDY4ACI1DJxgMguB22gDGZ1uXVW0OT1yYfNcAdW3
WpCvLG64jHpQzpilAprlQdbsdaOBJYVkoaUYdqeIBsRIiZdZcMKAQcJapkrrTqTO
DhyQY9b0iL7/TO6uPLYqthf2Ohi1uqrC4wsUemMPmmRXpZ7gz4sqzf6Qx3ikaqwy
GnVlK00X8bjhGfMtxz3Bqrbgs15Ek5eqA8foV3Yu5fGZoD9jpga1jyTUATBP0evo
JDjmbx2JzS2VhrqTG/45YeSHSBiZZX62qYvIJs64B3RGMS0HogL0D4M2xHfviYLE
+TU1bzLaEkWc/SIzoqSAHYmM3AiwnS1LSPajsV8/2xUHZT/MFtnSfbiIX4J7PzEb
vaVEdFbmVT3ig0VA6iQxGDzyGJnyiNpSJRxgBTIGp0Kn3wsLCCVxv9yMrRhG8s2x
a6l/wpZWnbmWE/7tpEWNyWYC9iTIkwEMdTICZ51ZUCz8bHmmmzY3MnHhdwsQLyva
MpiSQwVGHBRR3ccRGY2REyUqedGspuEC+RcWSZ5MwFQQPZO/eI+BzSDRCw7SwQkR
fjtve7l9VB2wX33NhdZpdvWAj0TGOcil6320SU9kvSZSuyJQLD0D3ce+iKvbp6O4
EWP/i+JWyx9N3vnBCtWY8D5Y31z3QwW43Nvq8OPWYd+rBA2EU/OllfK2wyVNRh4w
9uDG2Rrqhw8iQrsEmEjUZuXFdQGT4uvMBF3JK9Zs3d9YuCGfqLchG1D9ASk4RltL
S/J2jtFVNYlyHUyQUkkJg3FxiNamvB9f208Znpz23yFUouvTK6qy2mfO9CWKRIsI
HfmxlPh21KpsrcaeZbpNFUejky/gCQ7ymytd8FfT3/NUMFDgWMVHzZ10OlEs1a6Q
5/7tkUkIbEMp39kOSn9CFrBECGISRqkeD3+R/fgJek7in8YLRWnSGnKw9CsWoTAc
adhw78Wx6T0YBiOxv9/AT//wiB8XulLN9tK4U0nYe3lwJPvucMpobgsXU9aWy1bN
FJXaeGssYcI7DsmzV5t12JskAMepJEgG1WXafdcshOB2e/LbAwseQLlVdxp+mPc5
e8Rrfc7Fmk5YVjz4JReq9Wiw5tSeTG4vuY+Xw2zlRGXvVbQFBDNpg1mzrvJHJ/yJ
hpIQa5w4ioKp+DtQfKtnYinOY9F+P36EIGmcPm4YD/YxFgGc8fJbViNQ9ZcIwlZm
KjLDH4ybMbaC7ahutVOL0hEaLwZL7GdctIz4Q1+dfxCE3zImAjsV2fywmmdtrFyV
jmP7dtg1lGBa4/HshenWrjXzt0RpnZSRfu6G784hRWLaASb0jKvlEKtNUNONTvZK
Wb8GwZRqTatqsn5igLRwBEQm+ZklnLz2xQP9BZYrNzo+eWauKSq0Pwc/hUf049fU
Ex8X8ErkaJbUtTb7IMR5RNPl4cuMaViK7d0UHzup3YGJrjbrJE7EDxQcUJ6LpQvB
3GbqQqKr3EzqDA2U/q7V6ORmpmzIVgm871qIEg50q8ijeqibnFCw8VnntFzvwS+8
gjcNlhoTvSsEucBe+BsWobZbB/lJGg/EZh8vQpQvt9ZdtgmJ5i0WY3mT0uP7xivU
ea9VrStePtbQcOkbj1tKRRfs35rUYH1LOhbp3yHEOR/hQ7hQ0dB04L3+EudKVnBt
bN7FHk/nWiNPziW9umQTc6ZMOBlaE4pBjF7pL6bqSDLompaTNYWwegpXthwYLxLk
+dfDjfcbNFwdQXJ5J0kvdrrz42CPq7K2qWnskDsbM2M/qRKiDfk32X7zDUDK+qpO
PKAgQUW9nE0Y16iNxfP1U4KtOwUmR7drixZCniOZkqIw5kVXXVRlAxoREN+jOZFS
7rcSprj4yJrn781QsXBJm/E27HB9ilAsMk1Vfapfdnrc0xfIyNhYyA0zswmvL4Q0
WFwrBNI3hNJnZ50EnHIOEA2ISY1FeVvdhrXUztpPSdD4XxztUPL3UJbUaj2i3O1X
8hXPAdOX7UKoFovk4IrNx5Fuv9q/4hdlYMBS6h9gTw9bYSq4w/3j3x9YpHKqhEFN
tNHUY0gJQs9mC4MrmCXc4sqNqf6PMGqubGLtlKlYqmv3xlWbyMmRJkuAXVqIDTm+
Z4h/khenDQ8naSMZGRDGc8RYht5P8i08qRZk4AVLhQl0A+APO/VEI4CF4G+aKPoP
y8yMPwQxjBbB4kH9iDOfvH4EZayT+mm1TC8E0POLECOzLQ8aFrxt+ehqzfjkOU8J
fRWWt9I1Tp3q8d1F2cvu7BKV3QtmsIheE82EVzejbc+u+QmBDVcTEfbcjC5jvLT+
G5pbtQThxb5k0BgNKCnrLj06w/XRX06tf4y2ZxA6Hxi2gGzCBW8Gz9DGLiPh/ioD
572zE+TCr7AJXML4wuENah/v7AXWP3sV7FpDdXizAUXnxm/dyk1AH0/lof80ipBO
CQSL9Hee5Y0j+2sTLsUSvKpUaMg6VSsGHcipf6NGCIK+ABPcsYGcymihWaNllJov
jljV8GV0bhAgIfA4N6sexY+thWU2uBSRYunwTLHG4uELLKuA7nkrelYJZyd+UcWJ
haKOpvhSOgo69CzCroQWn6ymYXNn+WWZlbXVWZczETgosNX+4VOQUIVr6KyrRyVL
LWnZItNAcv/mgO4tsF2Ufrx248gyrEHM/9SAECae49yfEvdTj28QTRETr7VlHuwz
VqcJRj42eI1usXgfrJ4uDd+licameNZWSmuY2YFXn2H/g42kNoRIG/Ie0TaWw/ZJ
FCq9rbrPufO0dFZ88euLCi/JrjWRkRIjIT0KXlQ0JPVLMeaqghhhCEPUWOcnlzrU
4F1UmXCzEMFgGd1byk4HQNBeJsWmZwwzvAYBEwRQoEEsv+2REEyTwghb6AHO2M9j
molgd9WN7XC1nqizoPmwp08iaAp0kIopSF00/3GfTH4hoq1pJUM0UQBHn27t0JM/
yN/P+fAddP5IQ5/35iMloErGHLXhFV8TUXz1l38vky18Mzi6VXlVnK1F9eE95vDo
MhA41IAR0k7jBZzes7VzzOFNWkPYbt35E6G4BRBHmI9SgQQkaqq1XLFL+cBvnhsW
ShFiy714qFcyefcKUF5mnbQy6LbEvkNNfnc/sQ5DleCQ9JZBpN1kCmXagM39LWx5
ypD1Erx+dQn/OKSewPt+FUl4roofyHs1k10w4g/IOMCHxPRC6X/+1axG0SiH+iJA
/Hdg7tw7kC+E17N5qi2rQzvk0WIm0vbyEvU2/43KoSwmJLEzFKr55lcLzaAL3qE2
SzgVGkHCkAeCcmoGrUt/v0+JVxlQ7HqeHPt7K9/PKM4rKt+WsCIRqZRWt6K2r5Mw
/rMBaWm6cEdM/PtrqtR2KUlJ+TsecJHJ5oCEpI4ZFpwr1Z51O5XCyxsyZJQIzS51
LZ/ooMJdSs6ykeCKUfGZAVtP3G9eGw4uxOMdRUVfMbmY6PM16o5A+pVvcCIFAyY4
PITdy/HS3Ehd9S1JHWmP/HzUu6EivDzy1H8wi+0GP1JRqpQ9vxH8vH4OPi1b/w7a
5t7t9370zPabNj3CnyXaJiM5S5dD5sEebJ9ObIs3kbTGNQRbWBIEjcF87eqFWAGc
JPzFtDn5USxW0gwYbPKZyQgzXmPi6xV+nVNV6ie9EgA5yJ6CO3BUYQ5HQBGq3pnj
DAXA819cQWM25NyBlYjbwlpyIjCobD7wTV1OnKpuBxylutGXKPGsneogM2YFaeTe
TawzhAte9OBffHWZ/iDgTp164WYbKjCspcRFvKOVYHvD5/7xloiNJyYVj6VPk8E/
59nF751rSufkLU7gKNc9RGqohdq8tpvoN8tIln/zUOp5tcekh1E9dg+uH6klgx8r
QZ7qRFnIdFceVB4YTxHsIluw457K/2CzoJ1XVegXckQuK4ljqahQGoEQ5yw39X76
/mpCoo+T8LRYSLdxoRtEh2V0UJln4sDIrbQ5s27WO0h8MxKqX8Qx0CFXHvFpIES/
zoWfi/eiEwwkq72fEYebHCvlBGXOM9vadcMkwxUdqHCfxXTY12KIf5ZVWIxstHzF
mn8nwLNjuHc3kVxkkVvv0ZEyanXAsn4DO/zXVRZKdW4svVcoI6w4yh+156lrR/8q
ZQKyxFaOE9GuK0myPWTsrFq8g3Ld2tI+0uxV71rr1nzhyvXSbiWmSor5AV6/92p3
OhkWl0GkLOibsSg5+ZG41Oo6SUVFerawvYN1gd+hGlj1jszNzDcHwSmGy7HW0VKD
BmEB4itSwmS8FobHlIGTRAYeP319xJ5iqVr/71HCS83inusv3+1BNvTqsGdiFHDD
81CKCNVhD+3V9FZqdeN0aa1s6CkZTRWzbJyJY7NaMuOPtqIJVr6gZDEBwux0BFAf
AgfeGIec9Du+lclLQQu6RsFEjTJQo3hBe8PJA/ivCcRiERFi5AqmLN/mwg42OrWD
OmhwGx+gDBLvc4fK4Rtfw6G+M2qeehSE8OkjfOZlu1WnH+Ra1dS3ii+rw3QTLfOE
3ZCUlQyxrSftHn/VJ1qVL6Yinperi4fwZ/5nVkU8PxW0+FbNbRs6pXOPP0JkCJhL
lffv9lV4QuvfOu+N6as5wnljGBGio1hBXJqbISTBPdQfPLsszYsPKydPGHING7zx
JQzyk7RhHB4MUS0ul2EVJ7daRIIyVlCHvTNASPvu3fKErP4UZgLGlqNMsBEf1ZwC
kPdiFpN7V+l1k0cTXLtV9e4L8Dc0IpLdT1H4O3RF21wJq4UnlOkY8pEcEGgLcOz/
2S/W436d8FGFVnNzvNVdKZoQwKwkmUJq6KO1UMcB9kmBVF4qw8+HuJ+cqgxRGpax
6CX2oOhpvq1MSXg4QBkVETA/Rhu04lDlNF40sZw2GP2WmyCC3BeW13xD017JIeDU
Rs9XcrCyqtjAuK+ltb9d1iDAfsWpOygnlUq6pgQZPpvjMmqcc0SoQxp//WoajuaW
cXVUkGE3AyKRKeRWWHYOcpm4CWkBKgC0YndHHduVqQujhPGlaD6mqeLMQeL5TyWI
phhc0MH+bDqYHwQxCpyoqAL/M0nM69dj8L5VHCnq8OsOcIm6pR7KqsclG3y8uFZo
3IPsrFc0CV/0AriqW7dzYfBTOl0vKdZX2RBm4uItRXeR4F+lG7kI3MxkTvwplfIA
ppspsTiLAGleC/Kwxopq5oE0sbUk5xy3PMsLG9NyTLguqeMd7gkadX4yoMh7Hn2g
MiLwSErIu4kH/5znOoN7uNzdikTy/n30tOgjWlm/VTPDJLghbYbmNliF1S4efbEO
EqVMxNCqClitzOKvyLdE/MjQJ/UWdVdc5A983q8C2AQfL7wkORXHOKzU9Des08NR
/dLla+Dqp0av3u4/YwieMgpPkvcE2IPkHZ+ybLzOH8S6kjWDzZXLPtlqX5w1c1QM
q+bM9m2wzEXKUG+od626SSaReq/GDhHBEyS9OYGdUxl75LZkfTMm6iGBNgFU4PQ7
5MhYYJcRopB0pPAE5PpI+4iAZtLuKxF+zl9aj4ZS7AKhBMeBl9xGkqGHUYWAVKWZ
b5xgHCO44yxLh5rqQKBmK5I8VVKBgKo6uHb14ZRlW8/WQLxnq0wK2qNMzMlbgZwn
GXBwkO9ekHwIVWLN+ETFAFou/5nwWMsyLjr0pUKrlkDPiU4PF0L6h8ioXrasliad
Ud28r6powHfspzhU64RSrDAnwZS7809SPugpIN2li3Fm9qVwOaYmOQ3Bkpt5VDH6
XbkW1LCv6fjcQQVM/BcSZ1llR5yn5ZBf3QgzTCRANZW6RBFkgcX6baPaS64nRH85
wceDRqHVbX0eo3Vq9jScgKKfna3DUuD+tG2cCUUPkk3Vh4Dl6M86ELlNlD0pGNvg
k56oFl8Cw/snCiIE7MYkvKdeNZIAmvEu2ycN1nTkg6oz125CY9eLTVNtVk8kBC80
s8cO0iPNhxJA5rR9LwRrHru9ewIxx5jdF1LeGvIMnwI/yjnZjJr/1+BgOGM5nzRf
X1v2C3UIlizdIXYu0s5uNzcjAEgJQzGCBf/15WCgWdX6nIwZbGvl4u2DT0abmp+P
a3V4DbZJhFGeDPw/3QLYdGHcbIvcVWmlbyVUDVxudhPnqSWqUWtvWCPe6u82AdLp
AObMnR2OR16fj5e70vn8LJWjNWcuQAZyQ50YJUuRHRShYN+70zGQSbfX9C1WpPDR
gvv/CENEcyV88q1vKczFc8Pevhve3uYdBZctWqvnWWNrhd3HQRE+xnOL15GTgWxk
9XLiXFbJdNenS18yF6ny0iT7gGUEX9InYA7z7eH30AYpxdNY933P6QA6wc/zmSFz
26tgCKwZi38Tm9sB834TQBKkKBh4P8ZkamyJRTG5s5DHRaMAaLO3s+vcFhM+9q7L
L/cDFl3LLzUi0JEoWKiqUGgh8GTk7xSS3mZ06ErLbL9keHB/5VcU7GVu7aeLgvuK
EF+gPzVWiQRQR31/eU4NVMcAGi/Fd/eYl+TNh+6dSOFOWJDuAXKgzBCR62f98ihZ
TADcLbgBJ2qs+1IlsV5pPbknXnaYv7ch19n+FGVqJDCUCI4eJ29NrVCeoZ8LL0r8
/sIF1jK4vEnt1lV1fg4G3wtIEKeopV6bK/51HxMITwInE1taZykWx97JN/C3aoNf
qePQ3BmFkDRzIMcHAeiCWSvzecbqKARqzyHK2REDrGXqZnd/Fo7f+XZkQhQV5QTU
x/AoA+oQJDdCtx2DTdczooxfZfWq7pGaxxNWeUgHvHPg/QGyw42xRBtzLpZXYR8b
Xtx7wk19Jj4eB2BZUzRHD094U6ZO+3E++ukhsTArsoCO746fLajYd070NPVO/ARx
NjbIyKMi2hjDzM1eSkE9+rzwZenNWthl0AWbq+KeAfrXt39cMNTA92ayMSZ8iVZS
zLgazOqgTzpTznqkLdgKfi1yuNnQzxPgzS7JyEIKTghYLIwQn8Po5cMrM3cCa+3K
Wy2JILK5aeZBtpawmtNrSjnlgKN8bJzXV0scrHRFOjjmJI4o9cDd9b+ctb0EFSi1
z2c2JYqjX+cI+2SItUf8tYAOlTwcqcCVYtWZr3rZ+m9tEr+LAoIFWr/WqGJC7d3v
5EDxXdb/hMvOFNziI0ufiucIR3/tWQfYN4PY5EQdAm8tsWgEmOwIY18hu8ec6B0+
bnSQ3g5pYuBKJHkzYqfjQh7wZ5XHsjk0E5mXOPhvdFVH9b1Q6kyggA6oRTIYfKA5
P1J5Q6EPy5CUxIMms81cnJYhz44Db0IGIiqlf/1shIy6Y9LUi+tojWXDBFDeSkYO
j5lfj+hv5xXUMcPlXFh0gpEMQDF23IaAiBdgmvOkxXXf5r/1tMAF42TxgKRuDeSc
nIsj707PemmjRGNeySg+/vRB0xl9MFntCo0dGS8taUJRy7SmB/+cVUGH/DZKtQr+
7e69UofE8u9VuDZ9lZSIzdK0SrbVqbyNX67TwhMgy6G4GLSFH0E7M5hviCQLQwdq
Hgic7Rkg+20IrJtncWdQGNLnspW5iq5IA0kv2PfT/yPzA7VImSKQ+OAAOqWDjAiT
D1SQJo2McC6jjtITQg+WYweLSpe7okYaVBc2WsMu8Kn/vp2OqEwzxNV6yqTH8305
tbK/9VngRgAOFBflj7PFJkJ61FLw8ZghVs1y96vTfcXIArTMIwhFKd2MZVVtb5HO
JUX5W6ynC6rQId/Hs+L1I6g5Bq6Iy0xBcx1G0umG6ClXSB+AjLg+0zcBnsqEq9yZ
tdBfwP/r1hA+xlT5OqaHWLxyVosnqPIY3KJ2X7uPcqrZghWEKe/syee2zBNFYbal
Qn5vbewT0j7XtC+K/9iNj4N76nHwS+DXgzz639W+ufM0+6/sOJRWPtn14AwUGwiN
hYBRlpNwdu8THDI/FiuaGWxSNF8IGsNpc/ia/lChVXU/pzUSgqR7XQe+5K2oREf5
ZTe9mbScEEjgYg8ImX/HEBOkf9Cjnk4WAZBwq1xZb3M=
`pragma protect end_protected
