-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
UO5Q7TIWUFXNCWOmR41Mwnuw7OXd7u5U9CeQUZtDDs7eAH2JQPni3oc5ltc3gVDP
OPm/z4JpLt56NZfKpN0kT7qLHvl22A83IsT3iReBVAOvQLOjqUpJz+hAUNppSXys
Vfi+N4PYwkmTVczriqZBavJ/SVeyq+jDWa7BCem0A2Q=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 8307)

`protect DATA_BLOCK
475TlLFVzOLGHShbH97IzlHDBxQhM3/amDPvt5pB/CMRQgJ6nVpKO83TW69Y9DAk
UV0D9JchvWxp39owUVR43Zf6mAwLsvAZZfEdDp+AoVMPlBuIyTJ04vReGj2xen+j
AT6if9NY5TYG1lRA++B93Q9RGW0MMEXCT3nC2q6Gd7bLcaS2R721Dtaufuo/I5Y7
RQA76a8Go8TUd0717g1KgOAByyYp6ozbfSR+6P5DvAX8WkaJ9aJFN2cCYCt6HY5/
beAq9Z+YxkEygFdW5OfQdTcHoCgDWZpoTC9F/FVwSmTzwX6YqdoP97jnXeBP8M2f
aVWYCPlUTwSEQWkmjQHEaU/KKbsJHwhn/CcvdsuOZKmAvNEUFSFji+MvyHtCVCm4
L9n4K9y9RJW1y4EezCVhzPCaFzV+afsf0hyKkw6vPGEwTopOMbG+0zzKIBf8RAhP
uqTrQpo8cJe49SG8yvFcgfiqZN/ZDZiRpLKKNqBZliRo3XQTVlEkguYqd1fexzaq
2UQGIHMK3e48RhvrpkhrNRQejkx/iQqKjhgtBphmw4IzLacf7f9ugm+BGLKf0SbW
r4mYcSLKjJU8aOHbHw8JxSFYvRr/RPlPAKUNZsVFWeI1oh0z0chgIQKtfXv10LdX
mO61GKvUDw7DbgkEXmzsWQGxZq/Z4UC/xTMf8fd/xEvcFOZNAEN5kHnY2Cbqrdkd
toHq6RCjs2PioAkeOIavCLSmRKEEqXW+dvq4rWmIrL0pMSf8A0uXja/b6zRa8u1g
g4gaHBXTqjwBXYl+JLs6GCTFzydWCB3qvOlLmZF1PurI17tjp04w2nLWIA4zOmYf
afAEhSM0Xaxj7DEj/C6Vasr26V7dEw8FeHEe7YLbJhTFBpu2nkAaSx+B5EgySZtf
P+PCcnmp4YKfxkaG12Um1SwYlcgY/bTJrGbr8F+Ube/EF9SVeO/Wf5rm7SKwEEAV
Gm5ZLKx6mJbvGWeVgUUccelhQ4qF7gV/MXrpsxuJhs907RM9E+wU39AkKWqmc8QE
3y/fkyaU4qEheUHvJe6B2+z4XrFemu4t+6JdwmDGBZ8QY98ZLZYa8TdBpnUctXgx
l6RdanCPu6t7bkjDQF++s0L2c9QRtXk0C71nIhAZ4/v7o93p1BwFXXqK4zlrcI2O
4K3MNatuuZbJClrE6W/ER6jDDcnjNz6rbzKabUbJIkethHM4WesThQpHU2yZyM4J
k1rYnGi82NO3RIyvrCon/8OeX2RqZtzeJtVcz/QVUgWeWLwEjTdPNk147qv3PsLD
/B+YL2Q5nFl8HJOWUFfFq6kM2mTFb+v/7c/cdGiHCHz3V3ny9UDGE7Hj7FTKFTOF
Iq4wdDC+5OLq73d6QHWiam6rwSnM8PTc/4nnS/qZExwkGObeHAj6LJiuwUtqav8t
cfeNoI31a/C+UXe4F9kndm/Gvyjs0smedx/i5cE6uK06MVrzO1p7N2CmcDZQoCd2
+5g6b9t/HiOV+ogwVyVxGt21dT5xdFoJ8mHeCvKsBQ5ZMSXJffGfrDeMNxsNPw+O
ib+SqNbf/NWcI4zQuOAys0UbfdiamhVRCbe0dkh/1XjUtH0/xkDh4m+ACQpArUDf
qNc0ChQ9I4sCnJQTifPx2Y2RGEoTYzayz8UB8M138Lj9Pz4cGuRLVxWKlSRdtfSN
77Q9NZzyfqsWRj8ATChYHjqsqm/0avcqOZAlfikgR/+fL8lu3yyA84XF6fYKvwsV
SEe02SjFQnHB1qo7rPpRgWKdFIA4Rbz4Tq4lDgzJ6+cqdi8OgPGqJWlRG6a7MqaV
Njq20xI83o0x5xDXqbQqTefMX+HaJRn4upRZi2qETTOT775NKn1dJlfTWL35fVeV
TzMlL45+X1bZhMsXd6rdSzHj29RYB+hkHJF+C+VEKLVeCROCk8n9ru6D8djmnNEO
HJzVnY7t7jqNfX8lB17UzdadF3sm4IygbOWv2jWcTOoGd79ACRYxaLolrmvGSUtC
Tl0vbQxqwprvi58MPzqwg4DrXmxbdzdbegO8lYLOAccM5F3la6hP9DtBlZzuIWL3
AcnzMtKhZzwVEQf9XEevKvwifdPRSBfP3EbfnZ6Lka4uH4rH0MIoAvndARx02ZRK
GvU1un3dqtU5pFwVcLNz7gibBrYAoLCU26eUBTrguIYcwRALiybdbw3qCZo/651Y
OQFwB4OeSJxccI+mnmte8YUmyuqR31Kp+gS2/50OJGKm43Nr06iPmlr94oVmNE9n
MzZ/G2ySORvLTukiajcsTv6n3XUX/9sx2HY5/yF2SPxWPnKW9/A2ZinG41u06jkj
DIWLe5Sg8ma0gL8I0qJWGzwT5SO16EHINnufZ+gKghQVH2AXkq7zRiDjQQ2yBiHy
5s+EdhCQQeOBw0HSnrsBMkeSCeasyRtL6GmNB84HonOcuIbed5azPtLlbjYsHgV8
7BdZCA0usAp5iPJH0pc8DB83przdwGTEG2SaJhdYeTZZ1Hx5b22DHAPVap/aEr1v
aXaCQZ4iuvrSuAOHp3mXHm3CD9nOG/mR03YRPI6eJMCDZ+FOKaRLPxcLrIvCFOzx
+X47XE8dizRsaTMMyjiymH71OPU+efJtHUupbKxhEdEzEufy7HNjmPnlPHUfRBOQ
TF1owzvhEg3xiMXtZedme/Zomr30zUgqPnQ+M45Ujii+24+6HqfVVuXHcn/1oV2l
lvtp7urem5idGq+PjCaT2gCLpG6hERaFb0ZeCo8kmsmWNBK9N16sXAn+PgPm+hWK
ZoFIEoBZcBPMeH9NTKd28znl5P76QL40KvnFd7BLeKArsA/cPdWCGU5st6r13IuZ
YcLvn5QDbNK9GW6dlK29zwtqjH1c7WOIA+EShvEoXvH6tZ7nJgquMBnz/9msqBuy
1RuI4Q+vJqPHYxdbuaf/3qrPag3hqwSMH0wcMLeFORGbY/mOGDTn6e60QuT7xxwp
rU3aiQppMotTNVKPr9MwQbY5l/TMo/3BvFmzwnWCNQY+UScgwg98DXHUFfp1mjB6
M5Sk0l1gkf7ac0fogODPNi5tMhyOTv7Mu6VWlBUcggw/PQFbFSLE7V15M0mjnpnA
9Y1gxzRFfcrK+cOIEr+CL2NtcQEHQ8V5u3BkoYEsydS7ZfgFmr5XYIm9EYDZsVIb
lRrHq/QDAdFjSsra0ln+aWNjXoG1BRHIRZx7/lJLNmMGnmLPx/h0vy/APhx68uKZ
UPkmooyEkzUmoVUqwA5ejyL+XtLzj5SXoTsPqezm1rdfh5ncTkgxNI6O8/UoCiEq
J0QGbqo3eG+etb9fqc33y1DZ7Jdg5Y+kWjLJf7Kzy3RIlcc6BihQ82f6M3lZaeZ5
kFZMQFPBU1PI/hE4FB8Ozwen1W0MiYyx6R534V9/P5hCC1jJBJTYmjKiHL9G+tAA
i7+66eaUhMHh/7qeO4k8b0muMlWICVg/qJ7hwh8u9Xo522DK7bsrIPovQirvZcqU
ahhOaJIAB2ZV194y6muaHQPH3jRSER/qE1PLKtK3F1EeqZk9cXH3ZunvD1LH77kR
N3ENvNWKsAt0bcAc/KcXIc1IvO4Md44Hr1IRgNxGM2d7P25Ek+vUPmRhluFbJjTz
7UrDxoQULm8Iis1VbMO+IxurTi6hV1mzSJLtRj3XDR6lEoDKdor5I2yOPS4jCqen
fq8C3DBudkzc+oyOQPRUMQoLhhMDgDo2NIsxGl9A1KSjGSzC8g8IOL0UqwRhfiWP
2jO4tLqWcJQ7FiNLsBQFPYeJEa5fqxaBU1Mdn3Q7/AJ3PqoBJhewHiIIDCsHboID
dEnbjQ4/nRftmU6JA7rPlLWxacqLh6h8bj5T2BywvCLw37bas7gUiKbqU96No5Oo
X5grbtXaym9FpHax3NZNhBFuzqDZQF9rj04tixbhhKqpkUWq41hOHfPynqsoOoGB
JW7loc9BNyelX8MPkZMaciNv0muFbGodtZYb7DfWdBkkLMTM+bVq4/9NsEU7yvts
NPWzevA/gBZLXpqG0Wp3UmF9rYol6LR+7C2eooNBQsB1xUd6kgu8sRMbOTzDvmYo
iE+Gmf+Hu0Lnz8KrgisX16m6iHv1xCTeKL67PMkvDf4O5WnJm3UmRCTAsmKURMu1
30/mWDbcQ1sSjgk6uI3n4Ab/dQYuM/UI1tH0GnqicU7ikWWPVJd8ydzEdCTIokHP
c+EQ/oXrU8YfVls048JAG3P3uSuV8V/9u62QiQdRXLWm6F8wV90lJQQ0tR7cYMbQ
B3OR+glhKq0zcVLczhBqNOXwQtq6zHQX4UgMyW87Nq5xgpZDVnggbqGjHyvCBx7L
LeuzpkciErBlo9Ui4Iyf2nUeMtneW0d+7i2uF/BA6pgCYgVvGtcrD0Y0Gm0koHId
INxaFVHdMtM7GbULD032bBv9o72dR1Elq1Me7CiAKmNoVqteIHjujmUVeKpelN8H
u7XnpEv6nt04017J3lcYDtosA6eDhm9pAQfq73vNDvh7RP1Qc+UMeXUUfqWgbfM5
/Vsv/HT+13EKUj8AyM6sRR8bk2Vd9H95iEP6eDyxK8I5PsJfMTO3EKmYMeh1RDYl
7epYO8qCqFqTnRMm9PgTo/XScSkmCIDDA20WQcEGfKkirAkJof3wpbnpM4WP9pt9
2FhsDCshKJVso0whxdE86CmTCo0k4Di+0oaFjAc7dtoSvLeg+3osmrwGRdcFD16C
J8Yhnslvars/JTG5C8fGpLs5esBm1XTQv+4OuKIhUEGZLkWFyGJqvaLP7+lHTPjh
QPOhRXyJ9yCHQSFH1Ikz8T18amSP0rlGajQ+rBajdx29yL7t0rP00bPcdisPPrkv
+kYBg+r1FQRpimsX7I/lfEf3C6KSOdd9P27QZjKZs0JoPpa/Qt20ETju2c3y+xZw
HEZb4pQneVscGWc5WsHXPAAI/NTKCbw79VbCF/2zz10KCTepPHP5Ao7N+tcuNycV
yjOiMPBqHMUXfCTEhSBwtC0Fo7E321+xtQknDDi6bQUEkdVwr7b96/k5MFje3S+u
SlPsPMVXqlwraMu++O4ohPR6H9op3DnRo2uIC0YUorLrOtbWMr7vjSwsCuQkR8v8
VVWFGNZkCPuuubdqnLFwtD8smXW4s2XLSbHEpMYGn5PEkCZxGrc03FSdY797LVlY
OhDuMCZYkqpnQ4HyICzzHzGduA+diqpZ+PrtHLR68Vh3ru+NwMF2PkDDQyIsCJ8F
YpidxL/xug5dYQiBtfRheL+gNeYHF9vMAUac7z1sTZq+gEcY93QpHPIctz6m3r8+
1owd/gzDAtqSl1Gyy22M3bxAseMOixHFi4ao01WqqisUWCC6TCoNJX8zsj8wbE7A
SJdo8uJIw9MSAQt9Poj2GpTheW9Y9mFKWnL1EEAwAKMicpN5D+GDXjvSvZc6sZii
99UNpEoXk8lGNHQsowcMGN2A/1Y0MJ3POVY4/e8fMjMe8b6ceRs7q4X/Vs90wDrk
+EoS4CfU0IoqU6nxXKb+gGVyvgFk4GgvQSeH0BDth0b9gyIeci8Zm8H4evGQKYEP
38DNB6KQi8oAPgYTyQJ0GhBgm0efca7tqs6cuj1Lt2/G1gyRBYmXEOQTKg57ESLZ
zk9gzdq+vijYlqx/CUjz4klX7JL8JYlsVDPo1vXz8Q5WzNfCmRDp7dKbDCLYtWW9
N0621E4NK2KrfBFYoT0d7E6e96Od/bSCnSoICgpKJ5bIR14apJfr24SImGXBuf5d
u0T/VLoDpoTylmX8k6DggzskhIL9LBayPCWyMSyHzm55uEQkb5/aATQbS/zCtb1i
YCutjZRrsWixvSzbOYZH5p7Xdhc86+SKU/orPQtw0pH3qWjq7DC+rdTgofhwLSsb
5Ad2Xj41+liqoeXYVtWVc/NrYcAKORmXAk/Qg79StMuobBngUjTvQPazPOgB1z2V
rUboYYOFCt5H0bXYQHMo0FBudj5c8zQsussVzPE6vDdFgd9u2fXnbFWffl7pOy2c
jyK6y48ka3K7pNtLQ7fXClnPPhuS2J5XEFnZigb4nngj4M5L26mAsybRxQtGdASk
OzVIXSxLmejJrvmNLSEO28j2Al1tZESUprSIpgeD9RelKW2e3JqfG+K6gmEkt9p3
yFlp94wsLoakNjre/igZvizj4NY0hWwWsos0Hjwm30Iz2m/TL9q1P6XcXenyFt5k
FgmrQRnOx0UEkoabKupZnclYp0FCpudnW9DQP14lV+awp7BF+um5zT1OLa1/Hjly
nM5JzwHvq6M0GtlRua6r7r4TbwKnKckDxBHWbRebnGT7HMmXyOmy7qi6hO2yCSfS
0cuhRtgSgPhx0zUfcWVd4SKh60JP+eC5+Cfr1EKopMWHqfKBFaf6HG0Xs5wM36Q7
jQpmlv0fe9iXTMkglrliFxtGRoe7yqWem/P6ruSBheqVwAwFqddZ+1vb2bsoT77f
cERgO4JytsicSxGDlL80CpoRfjMMAP18cfiQMq9QXvHJyXkCtb/s7YxPGSEkJ1cg
6BhMKC1W2QNjqHkcWTfh0s7nHs8v93680ioOauAc8JNH6sAxuvuEN6Qi34+2oazV
Qo58dR2zzByiaIJVd7t6RDZmcEzwZZ/RGYW32k3vL3r6o0K9kPLQXYMf9biIA79C
Ufj7LXpSadq9QS0ZqFp5AseStCRgERyYxt/RObCDN6wtZqcMgDJ/6L88s6ZIYp/t
clRBM3mSsLwdeABRol9F+aPyy2UzeeQFSxP6gnodCeeeM9Q5wWKk7WljejmaeNGY
ILClROPokeSURvM4qxLy45rnLyYEgDu7z44d+Ytj8r65d+m5HY8/qM8vpAq/mjzq
xUYndThH0ydBkWHvvdZqSDHAx/XrbawAGbXDVE7eCbSPOLMPQs3NUr/qZ4NhOrng
NTIfhtwWcd7Iu9908Wkt6IuG3Kt8lw0jRTrSOM9Myv82Q9W8G6DfTa91D06Om4f0
VkQnZfUmBUv2m8xyPyx5godvwBcYJuGN/eYZPkkQgxwT+huPl8fybPXbr7pnFWaV
5mjVCrKrH3KtrxeeAo5u5CKH8NY1kvFTfuLqbH/uTKR/oWmRBSIZftKT37MqsNCV
5PpwasrFdwaVlHkIPKOtw3W7DwA7ELJ4xOBOIQP53Q2S2wRX2n44CKDhIG0qZeVg
7+SSzu8O6TmMcXdKldEdcoZ8yYWGn3x+Gux2na0LSqxp9hVra3HeY9Uu7x2oBT7I
sfLQYWHv6u2W4PA6h0dOOhkeRyVU6zVYMfLikvA7fDwjiXBDQgF7UzxtkDoQuv1k
RHATL6sx12FSJuQdZMrUjaX7c7hBT+CLRZ0u8/JwPQiLcuB0iThrgxvMNEKkPDML
xLZw68GovzxZaB6kO1zRnsauZeb3n+P8WXIrogE3BTBNhBedFH61RSd+0T6wjdY3
SAG+xBtKwg31OneXBkP/gyM45cDhailSkpuQrPnXc7XgKljdi+tLPxkYYxLFoRCS
GLT9sIGijuyMC8SpWv0h5IxCiNGnwL246grXT224bGd4Rp0NLRoFC1Q/uPkABXH6
7rF1U4C/LTGWVN9iOu6AKwIOGyt9ZC+YGuniOmFFNYV8bmaSEafYkvI9z3G4O5m/
QsxbHNB7dwSb3lgTMPWwcSj2IN7DCccVvAR9yDFPsID/4NP1qjt2sF6M27lhrFao
kQuCJMR57PnM25yo/T+nGo3dvJ4AH35Prg/dZvrhpQNErrpauHxka3Ypap77JXGR
rmaJwsx0IH0EYVcEHexkgR0W6araqXeKpKHP1CxiWbplYuFviEJXcN721oUbBGMA
t/0y9VtWl4Mcy08l7IYV+TyLSCDKEMUXqz9Vnp5A5fowd/wcvEXX3DMJeu939WRQ
4IXmCUBi2es52IIo/08W5Ep80i253JBxKE52DrRhlSq76ijrd2l+/EHGLghmaP6a
E0nCwDgpbigS7vVxUk0wfBc0WlNGzj1HXWDFTTECvCiInnMTTTuGQdtwQVABpk1Q
/tkozSKoOsFQa4pwGwpuZnBD1T6YqQTJOk6S1ho7zWtr7LmzqEW0EDO8rENX23sY
xuN1gCd9SA2+IFGY+Ybklhq+aT+3YvMJrQE1ZB6SDRuQOJxJE1P0KUrLpHlq420o
g479FXechPjgbO4i13IjF1Grb1uwLiJnX4uz2xANoxu6TWJ+05ivIe9VP8mxMyY1
6BmO4lbRfVso/Fx8JE6yxmvce7aDacYtdq0eGvSNoXbkqRaBZLbmoCOVROGjMHy4
yBsoeP/YE+cT7is4frpM7tQRcMSpAv5bWQnLhH5xaeesMG1QxYG0gLh1/20aNu/2
CNWngUmiXE1tCq7dgMHkMnxOqAy5MzjB1/npkVmStxHVXqYeg8EutYnpYuiViILt
iHZjq7rFR1inPJShKOoVHbC1zgFeSMJwuPbjCjZvJFDatfsiKO+cT3F+xWPrrE5+
ZuqNhSQu5+VW6SP2hdp1c47pWNkLsSE/gMxtOHD4OJP2g+17jLvloJjN27LM/CbH
Vl7+fwINKJLx+Y8If4YULN8NKK5pSRtnTwkNPs8P30FdY42Nhv94A9Qe4PQumBmV
n3Caj8irr4drJ7LGP5S5q+kMt4A32+JLrfNLk4r3qsxXbCpXzP3UAIY1vxsNMTpM
3R5rpj+iCf9qIdsoEfT/p4uJt9ZOGHbMaPWHI00SJSLvKj/o17Fl1+am3dNk+bOK
Q6FR1ar/FaJsmnkGBzMMpbAbWEayDlEzOTpHqh6Pq7szmsoPzXC8Ak7wl0Eq6ULC
kVp1JjLPxqeK22FbCAx718uykuMBVgHPbHRf5+U0nW263kUqjkIIs0yIgAVVW3h8
ijIrhSW9xpD01E++8722pWp3FhH63TKQWgH1FvZT+YL4dvYTOXF/1+UgCuWe3HrQ
va7orPyQ2woLnl6unmP82o4PncvburA4yybd9gZ8vYXsawo6HPcxpaf8SI3vO2Mk
133tppJ3UjobpWyiqOXqfQduZYnynAY/DvW56EK4O8/M3vMHn1MMB0HmaI7ZMph1
6XDluZaFW1DFSVjgEJteqUXaGGnFA/+PBbHILXmD58QPhHi3bkiR5clc+DRfboL5
igltJVMmJcqhZBwFfZZ17gh6WtwFiM6iU8JZy7KxYbnBip6UdR7jQ+vVcJh3WSAJ
hsAtoRI+gfYGkKDx7DGDkWyqNrw2EPUYlXdaXDLOcXBoarcQzqAIlZZR7ftx5/tx
n34N0+N6rq3wBRVRuIqq9MGDfBKaO/ar4M3KD8SnCk2WLC6pHVK+bkRF9XzD8cYY
QL2zEQoRVPq35tsKXFzkCJZaWYlvlYrz8XT3ipTXTGdyV93UzwUurH+82xjXJ+rm
tsbnBcRmMO4FM+HrjmuNVLNORLnWPRoavRQRPq/2qUxIvDX0FH4o0W74ExSuiDhH
74JPOx9Z2bcdKokEbrwvifB+As7Ctxme0cePCpdt+QE2MsVZCQcly9RQS2LJN944
BsL0GtDJi8gn/cpHQNcYbN11GM94Kq1PsanUpUYRJ3t7b27DsMdOIt6mkJyAXWcw
Qhpg+bAfd3KK71Ihi/FVnFNwwJGIk+qDgfCayZn2RMc8aSoXkeX+6LCSiuPxD05n
QmHdwnzQ5NP5blBOkdiLdYV+aoS07Y6RHomdiTuqZHzEXcKbdjw95lvnm432dGXk
iQXcUk393nCxiHaYrVBitra3YgH3kSsNOjDv8uxIyH8Zt+vTC58vIZ4UP2KasSa+
lgcRtRzKvsdYqtldVFgALCv5WHa1zZhXYRQ8hqCzFuNxD8SklTPi281nL+NNhmEg
hmE1SwpTHuMx9qbJ8Lcyho7edEg7K3gMZNtYGqBaTJ9RNHRl6MgKw1GG30saWQTh
hbJ9Yb0OApDFvL842YmZpQfoPZeCmB+jSjenMIYch7UtBBw/VlwZ4N5ameGV4M/o
BywtCpHaMyXWzhmJQpcHpEESJHfLOxGXx+wNKRwysr2dpNMvIwGT9XZFmmnfGlhs
QppyA6Cj2GdkE5GFlBw6BVafrZA0QLm6ivmXF2z63SfI07P/RYGkeEyY3ZW6JmjN
Q+k381L2ossRo1ReTKQsv7HkWI12HcSqmeHjyxzwKxI16zEXJKst5uvu7bV4N7Pn
j+dq3b5FLavSXIVKKYryb4I1G53bEXgqv2lEgdH5znmg7d6rqBFuayKVHYcAO4HS
/P8R/ciBV6ITe77FbGjKx2zQcU/ieh1NtccGfZ2l3NcTNaOhrYU+vm0Flrcg1Qav
VWWCJWnkdvTX/IJ4OM13KJ83tPp2OEf1IXo1lzICD/PwlmWmF5aXQ2eDN6vokUBo
Aha14QKgq4859iyLYcd6UMA2KP34GafIOiUc2vzN7w2o914Nb/rE/memd5SEy5ig
u9kIAoYqMpIxIv2cmtRj+qSutPYeUS66epiXEyY8Bfx8Z+smwRtZvx2NDqupW0gf
rO/XdJhiOAlNN/54hiq3FeokL0yggu3pA6/jDjEdxsbM2BC75PQHzCMlfmVyupuX
jI4RylkIsJLgb4sRZwXtwromLBD7U7r37kewvKD9OE7csFSeqi8BMEblI9Keq1nY
cbpdmwgRvM72P5GH5Fg6Tq/19S0Hzbl++l2rIoprJ7Ra8i67aXZaQ2JiWmaHeG4R
rx2en2TQzXt9zQXpKsiAG7Vs1uxHD0o4fDZLzGDI+Zv76b+zZEjIBg57TyYfYhXU
zrZYnxemEaW3zQGjVMOxRZLhgFO6/S1dlCAhV5RJsKjdo15KTcQaCSivf/HULhtg
fID+nhkklqVUxxtpuzrZnXyaqUIdh18rCmp5jQMy6Qrs9P4U+PKi3ww0vc812JBM
bjOnkl3QUUQhIjtOyGcAxVM0HdRv6bHaUOufeVkc5zfT6t9N2ecK3CCTVYyfXH0s
wNeRrV2zGz1LYOsHDNp3FpyQvXvTXNU0UyJ6UY6HH8SbJNvRcQ6BUUHqAQ2Xa2G9
iPerlG41mB1PpEcJgg8RF88m151JjPO2W29zIqoMSj9FurzZ1r2tBvsHRKjq5u9I
yQqiKrDEZXd7CmDrN5bHj/Twgo0F+tohLjMORF+eyOhkqqxB3JCvPPbdfIylrXZY
SSOvB07oGbTQsNjRr3mxjPWYn7yUjVm1qzNZ4bcUgPSY2wo0PwcfbS9lmjSWIAE8
WiflNGEA6vgSa6ZDI03/8y0PkYYWJB0U2xBL/RgYHrI=
`protect END_PROTECTED