// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Sun Sep 22 20:49:28 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jsWx7w2VN1J2ljojLTsJsvC7oEQVW8hHsgdMK443eL9X8rmGTFe0r1FNJZejSD6Z
1CWaAJgAYEG+BSksM74306RIw1wwpDeATEbusY9DQGKeCJm49vH8sT1C1ytS4dWV
jrLy2pnLrGq+qFUf00NX5P0yVAZf1VreJd2PtapWvK0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22240)
1oZQ64OtvKHdOKfsL9cNMN+lr9i9ymGyoZ+dBmy5BRi32tttdRrWxyuLqnIuKseG
zgRjJ+QxmNdG9jeCUh3eK0u8peNT5jvQxpWdbFvk/pQUahE+H4uODIVb30wk4Fty
vM2aDJFcuE/ULpUULFKi572x/KgZY5IIgWiexzelhh4qcZUxSn+VIg8mF3QTveWm
CM9NI2R9FRpJUyCTLPVhe1ZfPtCODeLzGJc9r8pGjJX+iKkZyu6tV3ySzLmTCVGq
Aif0guKWuvC0K/gJvdJKk2qoySzW7pwOVCUXBzPb8/6ShIEsR08+lPEkqh3jYctx
SiRhTBq2rYzyAcC+7jpLDAt1FAF6jN9MG2e+AfAdA2SGQ1WVLLYj0J+zuhdeE3i5
5tdHWvpAGuNID51RPTU3tewP3mVM1RWPXn5r5Em6Xmuy2gnKr23ec3HobxYBzpiL
OgUgKKiK2fSP3kew16ICofIRgWa1XlYum3IdauVu3PwcixQPiBBpy78oZ+kfHybt
IyDZnHgCk0L+1pSuExR4vpqg/BvLCfZIqZ6Fsw6/w0zciGPPyJi5dRtOqC+cg6oN
GiRwmfWQ2+rjG7kCQwZblSYap5gD62eay230O9lU7mymDd0Lq/1ecVYrVVCqA0WU
v2tlRfNPZBi6vkgmOhvtEcIeq0TmzQ7b66zQa95Q7pijOPpa4CIf+KDHHyS+hGWj
YqkE4kEMEIZsKlAnQIF/iXo+yKUasGRZU56XGgDCDrG/L802aIgvSpNskqQ18dgL
ywLsDXi2pxZ97YiACIwQpxkBzpKXEML4q7BNHbtcCAN/4X6Xl2puQpMMq1fLPaoU
qtMNRmn4FIKuzPyRD1Q1dmlMrKpVX5EmdBoKrgX7Ibk1Dfkma8w/UwEx43iHZC/s
UrD0ZNbrhFDvtoKnSTwsFrt5bSoCFA4oXMeTcgro2/iKODHUlFY2LRqNoW/BffXb
qBDodGKTXU8KOGla5lD7Oo65Fk/bd5HZFsvxoBiQcKfHAiYsTG+q2JE5EGRrWmac
9dEPm24m+wPbwe9d9uA7QInuW/wWj51Q0sWk6eGFLFfx76CFHibmgnGhAT4Id31Q
uyAKiKu9N9b92hQFmWoN5u0hX78zU2GWbMoACwaI3AoTk0cChImBug+GqX8zSC9C
3R+sG3Yp2QuU6t0mJ/F8e+rKodMleGIrhmu/48gwCPL93XbW58EZOprP5HqDFCmV
tEj0z2LQhuVnt7KIk93o5aa8U+yKbYr9bCH5uOWZtC+xZAgrlYPDYqUsaShcX8nA
USix6UL2T3wji4oahLujo0MhXez980dusR177WrlJ+yHfWlgd5WSB24i+CgcHr6L
RWAx55CyhVovtQ8ecr/4OHC6ba3nEQUtbVq5AnGRvhgaUbC1NpnyR273FSifWdfz
cTVKt/Bd2k+SH+d946ClpSGhV1fpvsoopxzqfDENNWEoQ1wQWwPhhRzDk9NRznyL
V6sTkf0FtMSzOhSJk0dq7QEiwoSUHFvtKDVAP2Em6f9KfvrJ1v3ZA7cfPrPOE/vT
FGtcMPjNkaaBvBPIYueeIQ676PQZPz6kjmDV72/WTZ218ht6wvNBoY81VqOqG9dp
4BGc76fE9/OAyd1U3L7/sz8za7k/jREotVLh4L9r2/I1rHILz7bbkZecR0ZnQUF3
qY9MDvfQaJeP2BHKn4bFnu9yk1If6o1Hv7VkX/obZJtt8GM1X2LwBhKySMKk878p
GZje5X30wM6BwBkBz4H5/ZJlr3RaWrGH8MVJ53qGtZI49sIQikAje5fSmttQmn5t
9IWzX8z2roVu2lOkkz8+l48hPlKDJGXiKuXdDZL3/ePY/0WsP7dxfdAboN2B4ZzF
e2bXWTxlyzbl5uo6zWaxwqpVDe39x/G+/tqO3HutJVM+dUPpEfgrWCbVaIQRtxxt
pWTNVTOdDIPmacJQXJNQir4iD0Sjwr6/LLkRTCAjnfBVjUw5zg0LWEEUWt4Whum6
BaIWxOPmMhcRtPtbPCbR6GC1hdukYgGhnENLgveYeqm6ziIy3EqQ6ry2msp2Iwf2
YRhDAVU5jtGzJJddkO8nXyAymZ/Tr4JS8TSHmS6FzPWKDa+v6pRk6Qd8TlcYfEtA
34VBHNg0ys5Dlp9Gf0oPUHyOHM7hpNa0fmp8/bcgDym06PaompsgANo+IjarqcMY
pb3k+R4sHeN6kO1yxfexvmqYRwnLKoUzLG23RCSjqBswxRgKGd/NYlCeFhU6VnNq
6B8NgakfNq0C2U1DuUictMHRy12yDem3LSZDlZhQGR1O+CmBpIlF5M6iWxRsxXN/
NTIBODcKUKD1wdJHBl2SkHfNS7WEWqbN7K3QGl85uoqdIbHw/rXYfJouAt+Pk+Fb
SHXJ6NqsOmO0DAvwKA1OIyF+XQTSUm/QDg+JVHFhk3aDtb1/OA4TGXB38d5zFSgm
FW6S8a3fqzE2B9ym3rjCqsLrLnuO1qQeqDB70VpzIrOIKecUmdHmZMQwz1KNd54Y
u3QhNErYOcyxFUDWO5hkKo20gYNxclZjYhOSoFzNnCGWOVND0w3LLQZNDwrGO4Jo
ouW9fjESx3D5qdtUEcRT5/Wcd/Zbk0hcHNlPvWB9vNivxxZsV8j+hX2oLoRp0XbZ
aG9n4+VQuMG3zQF5n3wUWEw/2deDFd4iRirI2mvouobH85ie5GeQ9DthuY5tQudH
nKENJL2BEYbZyb6s8HFr5GNKKzsKdHVyb6yptRhjCKV8JAf2PXZd/ARNFVaDKrga
VqyWvuRdpAyOW99lj9Jim6meU1V0FYYg1p2doGuyj/zzsFJaReSGJut+CqtkGLA6
yA3DoHfSPx4mD2RxKned70Bt309fAzlztOcin0CkGpaXHarouMzUFVm+hFCaotvm
16WhM+k6CVmmgoiVK7+KDc9hCro2o3Z0HlOrqbVKj6HLl3cryu8cCdHj4NIY2Qb4
oMMLVKhpICvW7+0QecSqtr7OP+O/BYyqlt6x1YjahwzcdHiWzsROm9ac2Uo+9/a/
l2fiFSVxqH/iD/tMs3fBKESBRXNh+jZIM1eG507er5jUk7aQCBdSIQamkiDciJWc
LFc9P3IYQPwTfqstcp2KCLQxbUnOtjRULHAvZJMiFPB3YLWsfK1yp+UX0G77WZkg
6/kuRe+Q/Qx3Af0Bwr/KGOZqgh8xoNcObzPN+siMVQZflvxE7xJMJgL7pKqm3jrY
gKqFQOoPCERMXbFgQbfujXLemeCw5WBFawjq3UoRz7kWhdBZIs0mEys/zxfIR377
XWPz3oF/Ls54QUuOgBqwhiHchHLimEgMPE7XMqwRHklUVBNPj+SSk7yxo/JkaAfM
/iW2XJ1b0KFv8kMhrJ+q2naXz4qNZjijy5bBzKmxUW/qbttGXwvMG6Pgx8wGgtxg
c6vLMPIbEOtYTJ6tJB9a0x3wz8+RRExaWrLqEF3Y4kQcc98/0vWhOEl1EQRN8SGq
P1V7IBvp3uDJT+N8uBF1sFhlCGjUdpZrgSQHv2SUzuApMF6LwiXlmAT23iY3d9wn
On099ej53qePnn4bm8zJUqD6STW2rQkqwjSgvzfC/Q0K4d6LIbC2PrCKvqDFbp8R
zh7F9bRNPnPRd9nvQqtnDrqzK++OoLafdcno+3WpPYkCwkReW2PKR+fI80qb6RK9
SFU++vV46W7VCw/69iZhkyiN1m9TfeooWf8miW7LsCb6PZUA1WFxcTmnaQZUKx9Z
Ws0RrlVPBWbf+J/1Nw7kOEF8CCVAuXJjYfilrHCMG9rK/OXKinzUO/jragbBUixO
saFZhjFoaVhsDkbgfwVBikAXytcTYHAZRbmsurkqHetdcQpGqKYtv0NcpEz7Zloq
hxU6uVcwvRx6yEIwRgNGTzbi1caVPfUJ5zE/6WrvPK6+Dhm8DP6+9V8c+nOZS4u7
0DfE7mVh+2WPjWq+Yu2r1YSzwy5RGkg9IRq90KGkeXFz33C/zaloFwxGf0wxleUB
qtdlcgWpfOrevfCR8v3ass+RS0zyrFmdKmJmEmC6lQXlL7cmSMhM6sJWGeEgEZqx
iilBf9Sr6QNHNruTgPURkvFN20ZlQvtf3wDtULsVokCnN24YKd7CS8GkHtScfWds
7NMJrVHCE2DbGvfoVDsHWh3AjD1STllNVEMv17DqsyIGT6zalyMAhyqyd3Tsfhwg
py3J69LPhTxJ7c4rTwsdBulXWm9fXgru1vR9Xftq3CPMFhL9/dqnux+jkQyF1PO6
FXBvTDpewdbyHEQ4oBvfK7rJEecoqNnCL+nTJA8BzyENWjk5z81ztg0g0cSW0XXR
TXBhagiRwBLiyqKSsjYPpKrvTTSkEl1F4gDREwsNpMlRISTzbiBpWr1xaDsardGC
iscwI10OPy7cbWJfhZSWVxA+fcV1Lb48kkvJWfq9CP16Z2/Nzx4ePlJ9Xfw3atAd
M54YVB7PLOEuAJPGVwRzrO6W3NBy7pWVeUdOAvqfnX84wpRFbTa5odUPAHqyrXIz
060DQj5nvM6Wvomzc80EWDfHt8KCrodcxmrLK3Sf26aelkaTkE3xwfCodRMuzMa+
Cp6hCf6igF3P38rHBCDNYdMj0mCiZZlPxINEB4yEiFDbwKrFikH/HySskMIhz11Q
Z3YN0U/21nBqaZcvKSM9QYIZ1YcyF14Ht8QLDxWYX2IUGS72rKU0PaHIGluSrF8i
0ClRknTPsazRVVOp2wFPaZvt4GlLR9ZxspKS3dFy5hP9wlZ/LqDYGhD0X1VwF5ng
ewOnHLiI8/8453XA2o9M7rN2qdwQbLb7rjpWUvF5VLKb51wbTYYAKwDhDzREAi6j
VnBbCjuUERmucHPFVi82YVeR+oBJwXx4rWzVzPWlmntCHL934K7qXocblHfc1fRr
tzk9Ifnef1im8utOYeXX7rdBb2ahDIzjYaheXkomeEe9qNN7i0nX/bEBvQSiufEN
P/R41lV6S/f7MN3pZmLi3mhrnsmLlhkDuJ6qw+4d5R2nJQilnSGVbipP+u4OTnob
M9hlSvpZP9FZbpYASvAskyv7iLflDIPQJnsJA5Ojhc+f2HxS7GZzGjtIoLBJisji
S0v2RJPF5O7RIyTrHLLFtpvEqYcVSdrLtYSJQ4dC++EnH1B3ubrqXzfw7DzdMBBi
wTSO4UF1cyAu6FOwnpAHqeaFx4q1iUGMvh8j/dOXcUVvxi6EFGYPpZ+60duBx6+3
XKDGlqu7mJOIZkuxLZzrdgpxBTU11IbJUun1qKNhulNGOGuUCKZ1OuP3xpmZ8LC5
ZfzmXGFnsiYYH/YPs2stmiJnq0oJmtaJ+oFU5MkF4CrKThCcbXPUzPEFIs3E7TMn
81Uw7ceqCe8TnzJClK9gpEAmIaS2Yc+pahsgAOEuIMZV0XPRIbmmYwIjAPvy/4x8
cfVK1Ev5SIAYE+TS4TA5dCpz9tdkdYTF3aQmOJfGDyRnw1vjiXRlzoBOyBEx19LF
wrxCOz8YljXQWwIw2cnknUEwNh/pVCn6PqsbjrGfF9yImuafJeXHI55s8dUNRp0J
v+y3FTs5V2L3M7fRM5WcQeCGKuB3gqYIx/aMFgAGFmr6uslW4jmgYUrNltJmIq+e
qsWHeI2O71Oco0vJhr5foR99PbTV0ouzwwNxXl65mc2MmsHmaOojxNbJ29HZ2s+k
sEkoIq43m15We9h0WEL0i7eEhe7oUi2Nj36XYQNR5/15fwMsuhbvg4RZL1bdIXSO
UXa5mt9zbxzEriHPkNL4IF0/vlckdea+mkoXGw9Nf14X8cEhVjyOAt8Xzv2yi6/P
VN1Xy6zf8Zk3tlQlXoXpa3Q2RFIHgB85x7QhkI7mvX8mGxBwW+XHvXNergZvUMgy
aFIzHIs3eQhkpnZ/uhHym2qHPrJc/9cYALk6qkIbLTKwF60tmseF08K0lKj1mRJ0
IfNruwfyRTuyCcminF9WQy4sjs3Y20m0hJve5qKb6+RUQAJ4iVnBG4fKDor32E4g
AYUi7Y6t1w/CbJJibGIqb0OKiVP7pxFWj7ri9Jvtmn09IS7IKSrMC9RhSU4t0GyF
Z9yShXOXNNF9ZfIEWx/HQvfbhcBtXVKhZKHodoBbGAb5Veec+CUMh63i7XO6cuQw
yRBYjxdG04ZmR3b8q2hxtnxNs8NXjEmZegk7iG44bBuIdiTm/Za2lcqJorXftINJ
4WIW+e2N7Le92PPu3b1i2e/1KwhXYwIhLdV5AnPShjBTLIH2WDAaiD8CuN7/sLLv
97UmVA8jPiUUf+P/l/rOVEIiQJYOJY3imW9gNVwlw+cWo53C/Fk/SFrinBtw+sWd
Bzt66CN8b4XrgOrBjZs65XB/WMmApiG+4gOKh53gjqD8nbGRRuyZBrHro9PHJ2IF
1SATuLNhmyU8Bevu4jwWXgBv7NGWdltRiqrUuzk9czJNjvR6l6609rvZTEoOPyhB
56d6nqPYct9sXs35+hF5VBuyU2JG9qChWqUOblATzzOw8evK69FeIVRJuRqifbQk
CAuDokZ72LTvqARG5ovB66eLYBVdrTdi/2JloByPcnLWsMw7mZRGX2S9PYXQjWTW
x6HmFdv6wePJ8TVzP09jL3/fuRqC9ye2vtfZjelJdwVhtKc4bnKUiFTlgoIi4nAU
qxk+1hyDTrwto1MEWNs08w03jM8zEAB9CNnmPDb4sE02Qo6R7Dk/VrQg3LBoai0o
+ExkozWLijRt+o3BjND19xvpPqqTLZxaWQ6vt2JjBg4+RPRQp0/cWhsX7ceoCcQX
9PG4hobFxVQn3N7BjbelI3ztV6mQYMOUg/lZPNnEkiHkNhPhiZKiHUBx+w2D41N6
fsdxaxgXbhcihm7XAtnx3CXTP5IbiiaMHkg3uRB1he00h8GEvEjQUGea6oMB0yTc
hC2NVv4n7duJMyv/+3c/pUkMFmFygDkjDKaO0fIWBzPHsPGYZ9jGpGnVenxa5MCc
uOXIF96DOEjK+R9QV7x1/24naKmmEShLTaJk0zOyJVNHD1oSa+pW9BokJuaUziyx
fjbKsKkNkOftLS3i87LwArZLkUYQqRRDo4YJMiS3wWUBucBtJgLeOTN1I0hEi4gh
S/nFdyrCcAz+IjPAnf7ruLozt/ElbHY2zBgXbkhGop9x8PUdDnR4ufJjDbWVzUz6
H+7yEXdJ9pe8BWB6LzYkBB3SpXDl+UVU00L7bJmyAKvJgjDEPoqxJyE8Q7cOdtUb
vpVs4/mmuCSh5K15Hky8MAeVvRf5P07rJ5uDVoOLUEEqqnOEfFCfzbcfNIG+zy0E
e0a1OJ31uwQMZNHnaxlh51Ta7vJ6qjC1ZpvuVmS9pYNfwha8gdHfMGuiIlDQCpLZ
bJElKKaOdGGbzGklRmPz8zXIbLmBv7u2ECnhpu82ZLPo4sshjJ6Q9Kp8DXnQhF5E
HIH5a4IO/wJceAS6Up6K0GmkQbapGZ78IHujjyQ30vmWeFF5mFfhD2wwTjsdHZhF
d3vw197AIWibyFJ+fX560oCGDbBjZ0jXzJSVN75sTHfZsehJl57sK0KHCUBIDVaF
pXnNj6P5eWcWuFvwfUnEz1/8noq/+FjYwzsJ+FfKp1flJK6pakRA5WemJxEFg78R
9JE/RyOSUEwAAB9hB/ln9m1waM3joswLpfVHGpYkEBaQjtWBwh394HgryhePA/nh
+StzP6qrM1T668asT68g1/mdOD8yrTXqgPEhXtLCvOBnnNhu5dLDAWPA3U70Zf/o
87mwvOqBJmx1+H/PicaIDnfg19zRUt+UY4L9vNhlkNQ3ozlDJpXQlv0iodwZNq3S
ZxcyxSMJWLo8dTcGD8zJV+IAxvOZz+DM2s2Os5QwFONIv8nJFv073thRvxENctKc
0J2eJJ3I9d35Fa+X8S7CV7IeibPfA5lXvFsYxSwxe/ZVH4o/bY8EQ4QbYgEpxWOT
/vpmLXDBFTCnrLrLmvcmOOK1cmY9ZPln9k4i2cNnGxJ6yCJIplHRSMpxBazCNG5v
m/yAg+fHvSqOT9plzIq1VeQQ4jeHr4Yu6iWdkbYwTm098Msgg4pw3v4LOAnLWEbb
hKfpKbzfIG3jbTkt2K6oSnSB0JBmQUUPaaUQ3JxMpui+BRKIRkEgpwvqEO6/acP0
92IvUhpkk8TSE10Xw6b0ABakAJoGA6nGRZwt1aaTbRboUbv5jnB35C1s8tKZIOjy
nq6VW7GMCvTWqixynAiGVfci+pRKvN7ET6RqJRVRk5AaxQC1aX2hSAf/kQDYhIKB
G9YTeUGw4q1/I0nRQkry08/NyJ7kmkNxX8XKNsiwJXidshDFwTnSvJWTGbSjaUZO
8BACqZEru8CXKA5ZYbC8R60JMyNG5fWPR/RZ+BhLAT1r7q76WenyQDo4INez7WcG
zbWJwVIiDTgJGpKouHhohPSv45mLEkbOaaqgRJwc90Ma5yccGnzgLxXIZVpRX6UR
r98F7IcE1OwNgZkl0rhvWpMt12RD8APmVKd25hXeODFdIoXSV2jHgsho9buvuFRr
0zXcnY+ngh3nzfEIhyfyXdI8bL0Ssq2yIJwxjdUUfOmD6uuL0x+8FBxSqeiauxqD
I7NMsbcBZng5q1dZlKrspebJ5QYwXEt9la2Ne0gplFX+JeqDYv5q7e+qcsLYE/pa
EjlZFBdOuBZMyyxe35Sp5eqRN7tzXCe/gBOz4aYnpPwaN1y0vk6n6KoINthZOhWI
7BYCJmfaIELIsPBiIutPFx/GcOliiEg2nhjxI31DWG6i+z472nCcZYxhla/IDwSU
qQvXk24rlSAdgaG/2X6afpfd7yNwSbODHsd1zUKhjPX9KbjV06qZMF3UGfzvDPv1
mOaQMMhneasowCZUefpHOqQDPC8LPLqAJxlC0w44ye0higZUpefd7PvXogwXof4e
NNm7kHSeLKngJKiv83KGGDzdJV6m4bCG2TV1URfGgERqVu9fAe5XDPfceNVmMDZx
WBzuHZy4BVLoBjJZoGO1leMk1wkGvOf/fNLSXYiO5BiHjpYs1UeLFyd4J2hhVuiO
Q8euAksv4FBOYhHBgVv6Nn+mcLxtXNK/Wr/CApaO5VFLZtRhKbIAUWOWLOi4EaBg
qcgfLXid2H+O2yOx0+/sQz3Otczdh5zQ3g3/eWCBcf31VkNPvIHpjymdMRN9PaKi
7BtxwaZv+PoDGf/CdMS8sJtmYuGaOk3d3jpXYuk5lU5Hwa3oMbOLFQjsYfDLvda3
+k+UKW+IfulmoaFe/tJpW7bAh/U9/MhI/k0Cb9mZg+SlEcEezCcnTgX9KD0/ep2y
H0tjVpOvoUVivIYRJQs2rgjsPZ5QGPVScBTvLR0ctZa9Ec4kaFK21Xf5/8PKEsPK
z+I5xBHmk91H6pqd9KwG4BNnKYn3i6KFY5p+fqQ2ljmtyr8A8/wDyXRvTZQ7xirg
RKXNkjHD0sFrSSFJrXkvSEBkravlq8K7BzIsy8bh2O+Wh1l3WmQYcGN/42GSjMLP
D2qEw+XbC/MNcz+b459Pd6uVDL4hFFvbsPQEUJAQXi1WfQ0tiig7iAoXmzGvTgeR
vjbJ+RkUDYCFvtcx+CDd/Yq4jKUbRNYf2yORIoQ6iDrOxl4b76FIqaz78iLIwWZt
Em5MAoptxqWQmbCWCKMXLFhK97syPpLFdy22ZYuMZHJXt5rXbNHOSX79KgLvSZXp
ceh2p6H4xgf3V+db2skZnJGwiFLm9RbTfn+Qmqqbzl1J/EuevPjPbGR5B9+nCeRm
PzsUJSRA2101s9vaV0ZN3zQUUid0P9mVXE8o9bWkzL5HMejX2DVPoE/HW5UO/Nf7
xIAsuDNsw5jKq53gkzFF2iuZ4mZfxGFNGeNDipKuGPemoIZkkWmKZwnCfTsyIwhC
Eof88JmQtoFkJQYmctI1m9LWN7UYnXOu0L4xEF+pyHWsXR4pSgmo7ih8CCWcxM+b
tNh+wKyDae279TykA1UAB6YlaB0WR0aQpcglCuuSRi5oICojarDpad54mNA+n1zg
yqOr+ns8aaz3K8qXec5jjZgTBYAvVfJCbMo9XDZrwmmLT9l+TSOUPVUwsSJQpmEa
yYxh+H9UW4kmNaYY+ZQKoL6axaR83/vzdFriHstpBNkTQwgU/o4tE5Bv7PIF8WFs
x37ewyyBIWK6thsyQWN7PoOPx7QtIOspfVjLr6dCTQl8yabcA6tUasworHY+c/38
6M8zIIl/kDlZ3xeETh8kbmqyfD1/OTXVEyS5cCV9kbJ9N6Lq63US7hhST/ZAc7i0
WAfCNxoIO/ng86Q4BEdqFbnIzF5u3tyb2NOGl/Cki7TvwOr6lfdBdUcTSzbx2zJ4
GanHN4U9Za6c0jjkht2uoSgi1PtzQa/kqh0vPeR7Vs7+pnh4PQJO+nNVipnYi2BU
iCPlc7qfBWFXdD/MFwvuLSmLu0iLRR2B2aLzTxisO1j6zMQZexDCIvN0f6ACfOnP
lJXXAWHugn70PBLUYBAl0p3REHCpIW4LX9L5pdz7+AbwTCgYGgtxHS+NFl8wyCMb
YYlzBjj8JyUzDNL3MxCCx1ukfx/PK58Cuvq9bm5FEugG094WoLAqRWSInZa91LGp
ynepHH+L1NsEphp16qMMsY5njNzXndHjGLZNUuZDn+WCR5tB3Lf2p//xjRoypeNd
O4SIv6fv0kazz31ufilrWOgXdE9RRxVAdmGlKH32w+Mi8cRFlH6wTanIhhOiFw8q
TBS0MUXSe4Z2vfs5vPYosGPn0q93yxuFhPejNC7WxJgTih/bNLq3w6hLWgYa0zAe
CKdsNdNFcbtNz7t0/otOYdDt9dRup0kF/Y0zNjKeJs3nTpX5Noh8GcH4kpRvXdSk
sl/C5zHavvb03NAqbiVsfMFcfZ/U1kNYtdXFzeEGqi42SSpxDSGAjhw1jd0TI/Ix
UTmrkUwSZxyTLre2PUElCO4zR6f+DXpwQE8Mw9Wbq2j0qGgWgpeXROKYRCXi0qc+
ptX4ASk3cg/VJ96erCnSOA0O3V7IumF7QSCDmyIcnTyWZrOaoCFWowk80tz+hSa9
H0ytMokuJKuE1L50ZNbikaoFcWJ3+yLbcKVe5P0Zemp0iFDCNw+bOm2Qgm+xT4cS
OJzUdVJKbpfWSU2wyfu+jj42kVDhZEeyeg9HHUuD+MumkdJ5NwkRUfVLEJt4t/fb
H0Ekq7/YJJygbKH6+2wxE8/1yPBF8y8uHgIjmFAx/J5UtT5/7T1m7/B9l4wIBmag
psBO41YAcvITL0D5t6vl/DO+/6mNj7oRLOGS4uAp4MxzGWyPN9FyfppWyseOljsT
ab07aU39yiUNOyn+tABCgElRGgmf2dYFTgaJvDcKAmR2a9kZgKO+1pi0kcE8X5FO
AxyB0UvWt2DAkBoYktqTi18o6+974EbWI3dXfvJNtvJh6RXB1wUCht5OapVIDlvZ
V1c9PsTcEp0snVSGtYLuF+0LaP9kBHOPTJ7VS3Jwo0x4Q8CM3VDCus9314YFPK3S
eK8AI1WYQUgbKKy7R9rTH9Y/kL9OG5q5afGdyNx9XqAHXWxTD8eiR1cAKVPeyoUb
Se1jNX3M0G7y0mRJAxaISirYnH217QXJHQfIIuIbesP8QaI2AM+N5JvKrvOaB7xX
Fy5W5izh3aWgGVrjfeVZXfR/Y8XzvMLSD2yANo2WabMnAgMFmXHUU26v/Rv7OTDR
OingtjS6mkPrmqhsxVWe1N9xN5e/Kj0+/DwcNkKT5F+CMH26rBB1swP1ybqTDlcV
38jRK3r3mhovrJLmHzHwvVabeVAeJf96RLpkZ50sf11bfpls+cWV23iXvP1DqPc0
cyvKgH5jQitLbD2geka2d5wYxmmbLz3X+JWywH+gvNA2fpDod6Am28pAtGpr3Y7B
R/A86R3iXSEou8jufV+Q75SaDv+3P2AmTldkbs37+x/5iVnvrs6XsvHR9jg8zr0a
lvk70FYeCKRuT7LMaYziePNwuf/B7tnyMMILKD9+A46PqG2q+5r4Yx2txJWaU9RS
n23G+8BXPy3l13GiwpHGrp04qhCqFvBbrF6MUEEzheVAAlAHXW0zNVK+opS1T0K0
GGiGDc6ndpw/8Xm0pS8FBi+jEweK3C+rdncb5tRiqQfkGECVJZsyq1BrHsMpdxI2
wOD9gtSO8HIBcv3+1GhtP/3UwmCVI2jLyo04wm7eeCNniSuwdNxLdhpBfh5Ldyep
4DDBjvvnue8/6L0GECruYCahjr7rH0PsitI8JxXekM6DZOjcOaHUcaSbFBcXDwLQ
JZzwAU4CZgY7vr36SzSsPcZ+llx4sSK7AM3qLmbFENefHy5A/kXRvHfy/NgoKFD/
qGPE96Jc1Sxa9W5cMasiCc2Jo+HWD298VzTBqYVhX6hZzQEvH4GAAUXjgkBHo0KH
Gsu9ekrh4fr/2XydIKAg474Q4P9voX14wZoEch/uPOJOslzXdBKVH0QDGkS/zlmF
ohN+drf1EqiOOm3O0grTNAJ6EHQDa21y4A/+4a6x8g5lfjSgjh9ZKG+SlbnL1qa+
eHR3LkmZU7L52ERnsSIN2ncaYHj9lKFRkYQZoM/NqtFtDJyrM7alK0ZDvBQaJu+T
v0diOVqbpA6FOOz+Ff1+gfg6TGA5hla72hi/TlF0kFcRtx3ojQbpoko0rpoBzJdm
XZHSBSudKjBmP1V5HFQxzjK9/yfrKEPs5b2zRL8zGd79L6Xd5gS1MPUsRElfXuRk
0HhgFaTqZjXcVSA8+kD+l3En3UO+WPuvrRL136QJchB1R9ixEY3kLlKHraLunsqg
MvvenAoxj3OIcfnHkc47ozfG5O5Gey37hpcuDSLoLph1ALMBnTSKQ81nKdb46tJt
8Cz2CB9KD0+UGLLGDhpmQ19+j2DmyTacrM3GGIZNYHQ43PqfSHUJJ50SoT8oY8xw
JieVxe+hl1GBvzRw4UBWmb67ki+C/qQ4cdj26SswP6jKDWcq9BjnZMJPwamqMLi1
bqs/AhWt/zdzKV7/b+7eZQ458Ws53EIIBRfOvqKINT6KNGc8Y2qRctjjOEcAuVuu
fHRkFNn6osbBAgaeDlla4R1BQz+msnws+Nskc9XfitwKQef9eaXPqgA5e9DeVA7q
ZgJT0CY+m1FBY+BcusVe66IkpuCXyppvs5ZmS4ai73GwPhxvKnfbSVU7Yv/oFdtu
eJwJtL6/wVABFQbjf3UmL9pr4TZ2MdM3oCDZRTi/M17vaRhsQxDgSToCaaa7G8/z
Cqv+0iyf32vr/4XrePkyFvIa8lfCF/p2ye/aYDbdfKfbOeM5kn/Hyi5IKQGJwho/
G/tk9gponpA9Zjmm7oD1aigbq7esb6C9SsU5fksBoLfQzGIr/Sh8mm5QXAH5WAO1
BHEhSqGIdZMiJijaws5ep768soq10YFreYi9gdnB6jyqObX/N1eYcyKkhRr/Vais
iTNXqKJHvqO+8NeCHhMurSobbHcDBdcILYsx8GzY9kWSy9gbjfyXQMPcOWb6EDLg
NqcH7XMT6dXqIBegt2X7Q0V52eA+tKChfgLcPFh4yye6zwOdsfHi/SpEj8mFsIXV
0NBniL453UQrPySEtf8q5JyYMMy8SMZ8fGgVegRAzTHglLF/CU6cbab88lEECeo6
fzqanswXW9OMfBL6O6AC36BZ73o7clmq/CZ/rqMDkA0spTPCA7TvoTn1g00THGNI
T/pSu843riW6NCP+rDAIu3+BGwkSGnapkQU759u+LjtUfh4ihraPVPEwdxbolqAu
Bngjl1uv5ZEI7RQ4We8o/WpgQssn00aVu308yD72VJshm6nOR4di1PfMsVSxnV/z
9GrqzkJnSh77MaoB1Et1uIRFnElD4HkOn+zsHFzJHCu3hVL/T5amwnMu2EnlCf4N
0nu5yOya0jmoMaJJ5yi8MPjtuppYPlN5J5bfnwgEApmhr7GQJSqi39r35l9q1NSM
0SKQ6GNVMfJnGh4t1XSHFIa/1sFaxSnN7dydvJXctmOaOyj8SUprkEZ8Ax27eJD/
Ay8dR0EmiEuddd0ksQ2IyulLx/gplHIeSJfgn5SzCxcQTM0NcgvPKB8/d4llUBJd
L8yEJqf0HBjvLQIU3W4J4gBngunE8vImyKDYGZQGWfmk9KoTtE8yvK24QRFIKlER
63Y7tL0rzsVBNj7cGUPI8xUvgkv06HXFhtVN6nPJud67QdmUW27r5wRnhNzWoXRb
Uhx2CodgaB6pr/fzIfDcDQPOOo8sQTjek5SQiKPscp24dUX++Cx8Jte8o3EWrwmb
IVfcRAcAdeL1dSmFlwD5M5OXKCaOh7xli2gZc5piPdOa2UGLycEDlOG0vpq3s6dM
bCeVb7f4GlK+do3EezAlSch5oPe+iFOnhZRQgAsLGwdDexVCWk+9Djq54iumqxJl
p+LZdNSmYG6RfH1ds9F/tuLSpn18Ahax9p2n81TWAYtt/Gm9zId5kFxZt5IR3u7m
eJJMmGynXb4ZdnW5/yllg5rymDLsMvFSjL+atwIEbXU+CrSRhkRGkMHH2absY6cL
i+/xlVHC3mmh5qEcK2PaV+ZdZz8JFuQoIOJ16esyjaGXQMaft1/8NafMxiT52415
FL9tmDyAzm4xgqTlMLdkeufpspRpeYov5vVLvIPglkPtCWIu6zKk51HkpQEhUBSX
5WE53hT6g/JA8McNd90MZKDF3Fy5cPegMD9dZS4umTu7BaAOnx5i1w/2SnQREJUG
Ot6csQiJRVObA/lNvW1qc533jRiVbmsPeTCM+rT1m86gFKi9qxH2giVYcSynYgx0
5vHWTHtdWIXzkVlb8p/UPUvvDD9EwBIU8wFqjBy9eUQO0ctYx1Bq1NjL+4R5Y1fC
XB8FijPCBiHCGO5dI35lYXe0WsfWD/6fidaVK5bhz3sJoYX8vlVxF1u0AJ+zESnv
PreYwxgm++l95t9lm7N9N6LmaXTgGucwwPRPoRUwYH6SzaJV/5CMp+6PAxBc0eZZ
e1VKG8zL0hd3bdnJVziGwhKDHBTNjIHhjwygM76H8uIaluBkiVfK/h3CXz2t7X4v
nZ/CbRcp1t301Yc+VQGHqHlktxF+BgZsyzj9Y2wkw8dmN2zPSIVYO7HvIV25rlK1
h9yTXIef4HUZcL2S81jG3tIkhcoiP+f3ofmEsfRdmBU/eEzLws4CluBRCfId5gXr
MFXY3tR5A3jtAE83k/grXT3iAGAo0P02daJHmQmMSOLLpG7AgXtmygt+0OGmhKbQ
ROrundeF8r+8FPgA+uR1tfcErM6osw4HfdLX/T4+0zX4qk+ZSGuIqSBONZCVuyWs
B7XywQeV9ebn/abcXx/sR7alWHwhTktLUbvPDG8URJdBs4B6yfMZ+Kx9HQlYk7dq
G3VUduQJhsUFDC4IfKv2pJxIqGF0Ky8Ounpg1ZvJ1TLQQ4kpwtnyL0e5DRO9/imP
4qguHzwVgjyWhfhkpwOCtPuQQi71UOr/c6VO17Z/qcfxcOJ8l4bBFQpDq4ITLrQB
LnmLfc0ZlB+JuCs237H0MdhPY57fmUDTxUyUs1JdFRmMsgpf0E1Ss6BU4DN7BeK4
CVZxfdZ0RG9DiZC4U9QtMUtL9v08ZjSQNjJRX8fHjvxM0yBIzb3p4KQRBrlL3SRK
pAuR5IKIry8XJ0pxomACF+n8il62udU2kk2CCbSTMrVkUZcGly25+4vwbJEamhq2
F1VQxF+OXW54pJ9Lma0LnePHD3BOS8eNOwM6q0wauTzYPxy7T8/gdwc5Dc3jaziN
pEKwmnM0S4KKZJ01j7SYchcbvsNfo5R5DH6vy3CCl2bte/8A/VgCW3hMsrSVaX5y
vXT1RVrqUni3pi5dK0AjZhzuXvOHb1e6H0aQOOCmStZNC8wR5p1z8fSGHck+r2aW
337PxMjI11swMdJ7swQvI+40NkrBaqay6sMsW2I17uC/7F5G6okhDoNeQveHQFGb
PDw1S/da39qYo6duhUlm1kqWeaVdyxgvyQvR5opBDGsUgUoYvDj6rQnxL7h+AN+9
xleki9wFJvViJJy0dFJU4iQHomNTapgAQzGVTUCj7mPIWroJVnKkcA2DGS2Tl+SY
bVPqhtUGinqq199draEQGeLQoOUDUIiWdeOSoh8t2DuL7wtfiV+2qrozBtzntwQ8
t9nRrdjFoVkyrEFssN8H4bPgXnn52R1COrih7/yUrLZvFPNQ84AQIg29utq4ouUH
YHMrRa7Ot5j5Riz8v6IW0svI9nCshCYAo5jC3vkx26MyXgzOLzf5uyV1WrE5opU+
j7m9OchJWe4ffFpYWPZ6/aVBdQ0HSL/U11P10gc2jnWuMFO19aRadJXFsSJvNCvq
mk0cW4kk1vS/iFIX2lcE6MKleEhq/RuFdP/698k0gRlMHMXeTjAwgxoh1LbA2m61
PvIVthUuP2BHgI93KkCPCNBBwRq0sbSf5IcM05g3yjH4o9hy7ZGXlH1ZMwPIW3jR
UieupzIQDjS4g5jMSmmrMpfrHuCOS0KitT+K9JJF58FhmwkzK9+FrQO1eG1zrJja
0n+J9UAdrvXV93XxrRRDpmvVnBNjUZYV4ozdIlvJ3KpoH1ez0U+o+/nBOd3aN9CP
JxHw3eB4skgKvZlwB4D6qGhRzhgYTC7R3SG0CmLUg6sX+JuVEOwoB/13W3JxmaZp
Qmq7ueFYL3cwzlFyq+yNbowkSIpy91lu6UTXCzZ/LxnTMFBbaaiGS0q16nr4+pf2
hmSylFMud7tzwcKwlBJLLpkdVI8RtAXIsGSZZj4afQkqpXqPNwlg8b4O3LlNJFdd
fuh2RcLqtIsFh4lds+av+0ZopsWD3i//T0FfBLpabwg50g+CCEDveFK3kmuBQhtc
pdk9qQFIHFXkI7jYIsPMn75JOFQOlAUkB0Cs4qX9aLuHqTiJc6erbRJFQVf4FkKH
S3Z9g+lz3duS2vXftbYsMl0+9AFyv9/x0R93QtIqbYqblLqq1nlqeyaRoPaBavSt
TuW4Wy2LBjwx3pPdVwg6a9eSflBwid+qNP5qidT6gQGckdMtZsGW7HUMTbPyDnO5
Ejx3Ybs9uFd9vgPcufhLTThAVDGsRYH7FMzBvb0JtgR3EmccJteQuI3eESYzEec0
UkeKpq/gfsMaP0fmo0YVKwjFnf+8S4TkZWJC/7dfi9krwPvkYRxBOCRBdKGtIqPn
kWCRcSZh6rQy4LmywyaLPcRc+sZAbCpc2HQacudK0fjEu23zjebizJdyouGgTvlN
W9hdP/YlgJjYY8acnz2Tm8SATzCaO6cpsRj7sylywfsr3qqANG4dsbY94U/moYjC
W/pWzNyDDTyNjal7maTvwXxPzVvyRnaLEdbUNrMNOwOMZXEWRubTr1kbOu0Ubz9+
yzhcyLnHD6ydz7UW8F2cjQDwBUKJDod+bJj+Z9MdyygSzAWNzZpqQLEdj7KD2eY2
2m4t1jHv3lvW7e46YOqM4rpU0n6Y0A0vTYkbbBfmS3KBVpaLl7x92PKXat5MnoRW
0TCxgfwwcosGgDi//huD+Gl24E4/A3WAaLCW6rtxgaeDAN/Kf4gXii2KJSdEvZRm
TssWQKqmwhGLRgYqHci8dHAf3QjFxr5HlfQF29eGQEs+Yxev9uJH2NAPCIBYrP2F
cMQuB90SJ/E9G9PizB84TFK+xCUszPi3nYj5Hk1RzFo+FLCJfXISu2BAT48wKXsS
VBWW6cnXvRz0XKs5JUgyFol0YmUyum8jwA9RPyiPebH6d7mz+a5oCbKhc3gbr6qY
QUoTCywJOHK4KiIE7kBH1cM3y2zYCX5FJ8CUTIb53oUShMY6RjnW13Ghuu/4T3Gc
jPevxgg9Wj2+wP6/3PmYtkNPYFx3WUanSQJlWT59a4cb9HSJnirvdUrOujmOVM6r
FFewsG+wKZyPRbDQeOwIZZ5X0reO1ppzB0BcQH5GWrwUeXw8w93g6xpJg5oq9H3c
mDo+JztEzKifFadjgsW8QUZpeUgSe/icFKj/hlrPUKmgfZ5coQNX/ZUsYSSAbt9c
nCEUAoVCb04JBqm2UO2gCy1kAcIB5CRxFYcONZ3lMhMplzqO/uUvbsZPoRYHFFPv
gfqZd1WdtjpaNd3dCXMnZli4M/pAxMbCFGh4cBR26doliHiktBQJtec0f299FCtZ
Ixy9ywQgmKZkmQJ55lmB/lvo4qHWwfGUVpAY3pB7Fhc/05BuEUjgLLtX8SStdWqt
cTkfIayDSWPBw0JRfYQY4xYuolg/JTQiEpc52/MiTO7MPmv0kE1+zY0uvRk+mmRM
yfYelZosYE/8nPJA4PToNsq5P1OXRf56u18lViwgmm/PlLiO/UxzRK/ltTvdrdHL
SBNthEjywoue/VWoUZFbWVyRJdjE5Y0JCHCqZcQZRNZOAQJpa9VedZmrpdLfAfWk
ZDaKqrc1CvGRGnOA1r8HnEpvBKnvtzpgV4lr0l5jzr84CHkD563XKaU0OrIzpIRe
J7Qu/f/gKJUUDlzRRumjP8T0n0YMtbDZyZODE+2RTrX/zr+IDte4L/jcKlXUS0PO
dO+lUQYOZKZioIBtTste1bCU9kK68S4PGinmW+N5rbPoVkF9VHUYg7RzYYWDWqZ3
bRBKDStWJn0gIAPoukRhRop073yBdw8pUYoszbXpcI2ohDchsgdiKC/QSDkmgNGU
Z1ZU3g4S2ZeVsUeDZ3YFlgAX1FuqK/o6Z9/6/QeGTDtXZSwrj3wW1sKx1bjszclm
Oz+Ii8jBS07ozPE18YNcoOMsE558Jjtgfo5O+GlXUwdaY6rAkdfe9SwcfVu6wqns
q+OUkWWRgOUi9hg9POYq+9/ze2FgowcECHILSySM2nr7uUyJQWVrhousTNBVo7x2
TPSzDFyGqHWDn74M9CBQaszI0XFfAmAwLzbDeMUiTbr4MXhYQfaOeIq4sbYGKPkh
oHeAt8pM2vYA6XD8iqvVQaLxPaYfMWnmcYUqkhLFjcVKJ7Z6JR760MBcIqHttFY3
5j2VJDjxh5/wBPQkpnPeqcKTEZw+rIrXT6ctRhhcTfYsTbTZef0pqoxNgaDySNvw
YMoPajsk8k9lLGW+KWhyANWillDEv4I3KyJnEjYtOJuDFhBvUxXZoJ7qgCexefv7
um33Xk0pO4UoF5Gj7sBxxYDpEe5hr0SRmAzzb96h/CNxy1SAsUu5z4/SkC6ok7rF
M4xAuBqlZFBwnTeZPp2NwEcxPLdD0qQvCxlSQeufukuJM+K6CrBYJ2IVJhHLq4GK
zDzfQ2tJ/UJ8fGA8iErfHaeXelmD+ep/OxJcGe2Rw3md47DXqK54YPXnhy7qpk8J
n2XtLPmdJBqSu4sW1QIe4kJi2y9iuoebZ51+TH77hSKxawbbcsZpUy9mEIXM/ycH
ItEmGB1g0caDrQ1P5yi3igSTsGz8bBJK7KaSxTv/VR+rPIZxF0BAausjJ/jSbdMW
0L5s/EGxZE7C7AhqDUz2gv8OKAhq1vbT8KcDlm+8bxu9Hx8/Oi+1ReDAaS2i/C/v
LgIeb0++zZAXUutVKAylBii6OVtQcIJlXjCwXLBMAL1Ho5lFbPSBQR11fpUQ30S5
FpNQAF1pQH7rC2LCzYVC6jFj5dkGQDdN/ipJBfKfDSeHcQcNR91iVsr++1HUfJ9c
L4gBueY5z460GbMpK+LVaLvqMzIbrHuCFEngBZW4L22iVhK7IXE+NL9bdoIVQnss
cM/z27LufBKLwAIWBqSEBB1VfMQKXHFVnq0UilwmO42dpS0T0YUPeJZCoxU/Y+BA
7NjOCzpDe7B24X1fk4rpLh9eTps7AVEKfUcToLPSnGVbQBSsUvHG6H2Qsd/2MZmW
n0THUuTV7axP+HTj2/6xAsRvvSvinYN+jQNguXmTLBfNqObtqLai+lT7DSPs/DjF
ug0u8GZmk46GtRxT2s19gSmb59H8U14UBYexJai11GsHDfjbadhrliCmgW8/sekq
GWDlSvXHy+iV4HRQLj+N4Q2cI5cYx2h+rlVRM7jFrggY7KK+FKXvH4PEYJfo8QCs
Pcm06S+V/dTyGWAC8za1cDAE6f36S/nPCKhD743TVRqZmfSx+rtZFVsV0mHXeWAn
QsxF/+o+R3/zVZPwXvkbIlzgSfH+QAxHSpqu+l2SL9AF5rtyFHjFPUY8VhXRHmL6
sWzurcWB9gNCufJSs5UhgFNkluVGS2i9Mdn6s1Z/kKaZWA4vqFXuNjcAIm+4I34E
RqkwYtN65bKnBWUNWtFvuepyaZLYUb3bnuD8SvduQDTN1ES9iY7WkPP3easY59nY
olA+bf+q1h5sp7o4nCfj6SW/HspOJQ+duneh5wMMe5fxp2RTqVUzf6rNNIIb0ByM
+SR46C1IYAE+VCe2SZbGmxFoVjFKAJYXfFlAl94jKMSjpxe+Kte7pbQyKdoWFrSl
/pCY+6o5NAAVMwpciBrlSJLWGoRAg8BkX/FbjjxdwZorXs0akByikGY3Ndg6+Gvt
XT+1BRGY2G6MOj3qRf4fELtfN+SyqmDost0BERe5NR/QMf+xvgOVYNcuQSFnG/C+
5ti0DrYcAoapDalrxiB12NvKWpWI19GufDOAJbvXayXasEWekK5wTynHh8QjzEaC
CUj34tXBRg1MaDSpXN8olndKAjV4WRnkYw68I9/Q87gJo3RAa1gD7GkJrHuuPpya
fP/G4vR4TRzYyMDD7JRrVsbHKPHwh+2GcHthQh2ql+wV0W5Y6jy7RwXNb+lowc4F
sjQ8uGltpSWj4WC3E5PRBuPSQKT5D9V5vKwE+R7Rs5Ptta18zx8XnOB/K8oZKHhH
st25EAAY8tbN4SDeBHamD1JQSY3q5HAWpUMCD3/lwbBuT/PVUfDNq3WSWq7x1gR1
QCXdKLRcEZWA4SohQlhI6NzYH1cNHllZ+WikoJHYMdQMLZA/g49yqOWIu6ZpKmHG
ZfPD5i7M2rnD4wXerbKxWtb1PM6IxNzFAifKmUwuDOeEXsXriKaaimdDqbEOJvsO
4LaLvhBl4Uqaw5JI4sW9nD7Nm3k4dX9hdE5WIXBjjMBZe0VuWkvxHQLhLx3egACP
+z9oTrokGIKNZb4ON+igt9caYBM6qfTpSFESI8jvgTI4/qfuwIZ0dCvdi0z8L2Ay
xgPGbjsBsGaCSLv4/WunGhW/ttfFlY0Dn51xJ/KiNIrlPWAadUjLCiTRYk2hWbnV
jnkapHRLhvYsHdo2L6R9lndMXaZ64D8VBsYJ2/dluXqkb5iIALoAyoxYK/nUzfDl
X/cLTMisULZiE432EHQW0b3gtJSW1cR+r03EJB39J3f2VfMafhVv+tlgtDq9Qae4
6unR4Bo5kt5NyQIXJ76R6vdlgKMwDoX+ZzB7OdD3Ev/glZ+CFfLdyLoncf0miR8t
p9N34tvasYY9GHBRXQCI2ok+EMssxKPxJik9evietIC26brY6ckZ77I9Ac4a9k53
Y2KhYhs4BUPx2U9SNqX3uN0eTi2jS0fxebAqEBsBHGotUOf+wssdlggXhpmJGbvd
68q7SyI7sAjoxKdtPAOHawigpHYzx24WhxsUZ4LGiE+yiMtO6d46XilM8pRJhM4i
lpDIWEr7UKN39JMCqb1tl9d8yatQp+e0lnHkDD/PtJ0enEMzc7eOlf6sFJVTNG+J
Q9XlFW12fhus3GnK68jv9WrCH9ZFZmtg72TsckX9vHUPsBN3BhLpYYR5mdHt9JfJ
45S8X21nAfPFVKuv+A7EM7h7IZkMRZLYxA7LYKxVD1hFhXV+mQUiKDCCUs7wSUQW
HEjovylsFOWkxFmtUCgerI++ls9/1mHW+amdkzpg4jPV8TwsV48EIBON+zd6ixt8
pSFZTnJPxJca2unOGd5tAmtgeuQBRWLP2eT+JWvNyfBv9r8S8iZWWgvux6SjsOZ8
brz94NLv/EeL6ksxj9cZm6sJltz3cEvl13p1semUnjURFYXDiIKGX6vq6IUtGXUg
p0ID2Xh8Wpk35qP+/xndu6HjhxLtjekLt/QIdS6xlzfo1hMIOcaEFw/h8WfiCJBX
RDWgijBh5GuHJrob5HtEI/l2nIS+TM83OS1rByweLdkHE4YJsHcR9M6HKtJp1DZv
I2wLcWBKyFyWki7xepvnjWrzYJGdNCEBeeEXvBWIs9boMT5iqUM+rw2L4HY5MEd5
bxCS8uB7m8KXZmgXAFoKhYvEmuT/UegTSX8W9b8Gos4wNp5ik6ofxEb0FWFgWVHJ
Eewo1F9wQX1RjyeBcDiJN9IBkFFQaiQJGcg2rdZGunn4n6kHY4xDsNiY1P8FYOfK
7fTYdYzrvaoEYEsgxCvkZg7loGQ9Yze7FeOQwWqr8GFBST3eAjnvNzBAsoUv7X0A
cjzNqejH2+jK2qTY2F9kScJrhxFPa7m+h8Glx7Qaod9vqpdZaUxJEtc4Bv2xlTqM
Ddb61QNhOFCIAZTiTZNGp8VKhRxzuqHUTAMg9gckTp/FP2ZGeHf//dOTZk6NAZLQ
Iycewi9FHVIfAZkbqYfJuQeABTYCyHn5gxYmq2gDJCnEOpMuT2vfj4ViA8joRe10
S+svYiYEcsD8ejtaVS/+/Vh8/cNb+RLUS7FOL0/3bMH+WhMjGTQ411RKpZn8TzQ2
RV4g53wKBb7ShRSCpcDiwhxTSwqBQRqyV6pijAo0MBEwF08whoYKtsdXpJkC14LM
bblJFE9aUgQtiyUWzHPFUgxVw810vCRL046oJLsQXPypyFxc6rtNJ32BIXYI47q1
2quIMcZTIy/k5XIwwCyrIcLE4Zt+A5s0OKaYALeaI7eDPm5J+3u4PJlqRgIudFT+
iquE5gD0njSieCLIgleGVY2njuZeMAsPzqUCqMD54V3SeF9dU65OV55eFRMJwDvu
Hmt4uWTY28FX5GV1dC2y0p/noc7NakpLLdrZhW7uKlVgPheqd6yoSylXPXctmc2v
DsSpmo4+QoPjIphzhshMWcYA3jnWYldIMGIVShV77N1vM5QeDb71TJvU3Ud0b5Z2
eDa3tsPm+sLMI91Sta4MrXR2LS2HYvtLukAkkhJkG25Jbtgq2iPyOqfHhJKHR2Pv
ijwGPcP2i0g2K3IRHe6TRVmfiopeUEJCyDZS9mhgmZ1hgPP/g0/+iO4UR5IuxJzw
Uc3ryP7Clzv0dijBVuzPjazWoAQJOjAc5vJ/wpLHTx6da2/0KVzITU5hSLKY+DxF
zfOvE3lBB0n5BzhPmOC46XSG4KU7mvC7slgrzuUcg9NhPv51suReoQLMNBy1k66o
mrSIOtaC2gkU6W0MSzIFUv6R0q8gfHdr2Zaz6exzNSoHped/x7z1dNIAhFsR/Yll
5ppBb8eZ8wdOQ2skJJaPVYCcOjcPKbngEKeepa//UfhHsNtxVOqHGSKEbk1x+GA9
ETeg1UBj4iXek1cHQrPz/t8mfYdVFemdB2HreaOi6N55NgxxBKZjO3GmBe3hnx+J
iU78lOTe2PG6QfCjNp1kSryYuvKkVbDayMVEsDt5mTNlOaxC6E3iThzXLFysXgvY
KkPFXXv1jDEbHg6PdJFlU0CxB7XQjR/mXTLKKi/6rZ9kKA/WXTmmw4mAZIrPUcct
cfPJYO03n7LDM60zmEG/bKv/VZX8IQ+9ASFcqb0lK9ajif9TAVKOx9wGaVCy17gv
Klcm2lhRQQX8YyHMXCJOaOt2warzqr01JxfO31dzUybRsa6NIQN4IcMHoJrfaj+L
GpJ4nXuJF5y03sVIWgiyqsINc7hHEs8TdNtZcjKm/peBjMRDPNqeIKOfZgl2FqCq
Ox4+wpVDqnwN0WAIdaz7xjbR9T050LtiTtn2eITGX36n214dmRyZGlZUP/jq9lhS
217FlYER+PlWDJ1n7vDz6hLPxmjtJgTVqBrK7PuqwDKFa5j9einrt9J43aIZ/8oA
bodu7a+e8EF+XRjE2FDL12DFjS9gGej0KPBsb/JZt6uSbOCZlsbxdteKMuqSaEVx
56CYBTbbsPj1at1mMleYKmJRNXYuCG2j6PHIXBWhal8682Va4XStpk/yxIUB8rpa
vS7vxUBKMnWnIyx2KKVCFtgF3dstELFZDh2bZcMfqBfOuC2vyNI60ekU99VeiTf1
qmJOZcTcRrcEJ4HPfmi3+RetLn8kPwFA7tyrg1RAXETjUiPwWnEA9Up2WnPjf/Bq
v0djINseH+Pe7P+4po0GSwDiMZILAhw2P/0T17XaIqeSdc0rrIv7xmZOq5Tkl5xi
npCAhlH95iRsI/eXUbjeEGDqAWKl+ev3HX8oXBBx2GUlF75nVKVzNND2cxWWhx54
ZddJEtC+3GiLpXQgtmYdDJjKfo/96Zzd3FVLZwOT38jFA7yB/vpu8P10799wM+Z6
xA9GNPjpkZt3o/bUWenz87HMvu5P9iQeP/iBysXzDQfJybMKbgZhXq2DJ3l2+6XE
TQPLvIGZEmcDOL4TSzZ89bHBrz8XsjkMb8Ejaq+pqLNqHzcE47bL/w21Bj6dkso2
xvfh4VV7ss9NWGGpRr3Zp15BiV9bPxvqFOodWnsK0TqlUonXwnRWGUJJ2JYOKq4T
Tt4id4SxVM4p49Ugap/DDerC5B7zEbVw2b9COagFecwtGnb3iyeL9C9Eg69qQhTK
ecxk2N857TBK+rZ6Tz4Yjnp1Y/p0NBTfFqK+g5OH1NYDSyefq97TQf1z1FV7dksq
mibsjCZKlyzwfo2TXnnsQrjUxZPv8a5PEVvEo8CmIgXnUrwG1luI8TCNILjPeoBr
rEJZ0iLg0gHnbwEOF1Czro3ml59gI9Sh+mWmTdnYJYoLavBmRE3KTWv+d+RkpfGd
6ZW+hbsAfTZJmbsV/PPGDYgHltxiRdTFpatyK4FIH+yGRRMCjzJam1Cx2zSZ1GA1
kewC1CAORd/MXhHbXMMI/tjv0yB7j+McNCgry5ME7BiL8dYl3DTjBUt8eg9H9q6g
38Cm3hRTaw0kDZXTX5tlbBpYSAnMdMz3nZYHrMUX7pHmlFTVXrqHnSUx5/P2XhI8
G3aPV5OHasKedDaZ7H8gd8QnCDhs+9VmpgPJL9zjWQ+xho8Vp19zccH4S3qzbWrz
92kci71JPR+zabCP0jQpRp1IXZf8cPZS5rzqLvLfIi8NnHwy8MwjK9xr1fuO5TU1
4JeD5S+GnfNz9lCdZtEVgk2mVs1NuGNNyVLnknxcyzHgQCpcOHpbZfncnDu0fHQY
j1K4B3+4wxbboxmeUveZFficZj8fgb8YGTxA1muJKCclG9EhrmFI4Fn9YooHvCzq
SGmV3D/NZ3sHCv/UZFX5VHnm9nBf2OVLMjLv4KsUVi1GVh4P8HoGfWwBPOA5Au5I
yZ+LrAd9ijNM9QQwWxKBKjZ5/NY4JBXizIqnQXFsFiJ1LNUFQQvzs2A4LtIxFxGg
rrqxy8RC2EVG0BixfctE7deK1WlL5fBXSaoeagB5beGSQcWdQ056fnn9Gasi+kSg
yWtViwvOpjU+j/lxGSu2WYBp4rfxafsBjlgQn+hnrC8uPoTXwdTilyXAAEgGiPUr
huO9BhBRqQYmt/Pd1BZhBr+i1MHarx97CWm3pCNWL272wA1t3WMoWELNe9C1NviY
O4vs8QVXbwiL9B50Pi/ipLtu12OYdcH2P9K5Yts5fKggyBG2ssbLcqVmq8dQwDzx
iKhof0AjNET0xihbAPQ3JOkBtQT3YzYIATxi6wCt7zn8YtR12GnyKMN3/S1JTiEO
4Fu1siRINubC60GBhFYjDvTx/rGPAHcn/XU9d/RLN50f7IdI0gspYp+LE+YGZWf6
0SjUaJJxU9yjSlt2AbBzU47F4Zy9r8lp3/fLAAZWoLd1942sBeZO7fElxU3IoZ/9
RbFSAwGewFo6WvXreG9kIY0PJmkKFRfYz8nF52nwRMJetmnNA8LasrUoTbGodEht
WJ7pnT1jZyncFHKWLZPgF/ptvA0UVoT9aXM73lLO4hcTUm0QuclIoietRKhQ8aE1
hfwYbTnL/6fBcFG4xay3GMTOOz9AyrmZu5lDjml4k3kOtXJDYzLl08PYH8ZdP+/m
GeTWns64SdjZxhoqtUTWQZf0mUmweFAa86EkUngQgdzNXXKcMUNXVk7V8iYBt47d
y41LCj090VzuVDgeOJhuZwJ1mWTe5tKBxzGQzYIJ19AC3gYdzjhfZFHox0GPfeHG
KonaGoZVldqEysHfz8qkBjqPT6Mq4u4HjpsIB9wKM1H3RrosuNKS8TA53VPJkKuf
kb0W+s/hKlUpiQq8ljtCWRMfacYxLMu5LOyFtyf6PLO6D4vOv2inCuO5yWqjjydg
Kh8VHW9BUuU2QOrXAiakJD5WD2Ll8biJbO2QAlE1rW/QpS38vbESiwnSHaV80rI+
s8EuTtI1NSH4ZVTvbW6V++5ACIbO/QWxB3vrkidqww3RIbM0+mmHZYDDmuYIYL1t
q8fyaQ71LkGnKdsGtxIM3PYQJH6mLmrhkGxkhCFW4klSLBsmrvOj7fx0lK/idOHm
cprEa6evB6eeDUC2TCbFud8c+Qpa40sfVZ36hX9ezYoUeGPCqHm31xSTL/7dFpY4
aw8R4WOT/xyTfr2wOv+exLQMeuqjRQvYpEXHbv0R5BBM39X3LkEAIPEi11dYnQFu
aKQbT0pPSnxe3ChyutteWTA2ZfwOUrEQq0ng+ixouU3UqgpKXdAF3duptArnIz06
Fbo8ELOw2Vx2hxBBcpDY/vDLuU50eCdwUgEoFg6zFUCaa8OITUVfVwTqIAnPtsr8
lhcCjPZ7uGaRbKYh3PBCYlf3NaIyrEe5zwwBU+ItQ/DrGP3h68Q8Awb8d3pA3O7P
SE0GvIN3bdcyb7tsQJiD01P7AtI0U2N0rddDWiwm2a/+fLeUT0VTsfyt86YbQpIu
+RT6A69pjfe4yM4NPi9o4GOY382yvgu1XZdA04Kmo7QEXWbCumB7WOdgAetwhNdD
uxIl96oZLBnqpOlPMBeJW6Innx6aKvTjl6VshRPdtj1C1Vofg+EXOK3VolFhanUY
cFkezkExB+Z7KtLNEDzIXM2s2uorOT3aKxYF2s6geIW069vannhdl/SAtLhWfslO
Vc7sGS/+tl7giZQxQ3wjReTkn3OrzeCCYAGzJoOfBCyK+0zGD2HqtnhCKjI9GwPM
b7xDM6wKJNXMvAYIQDZnsS63RUWzaBBYUWUGNJjXNvqRM0s0XzIm3Iu+xXk9Q/6i
FHph5On/jqPMCTAIsyfA0YalDvf9aoY0AvRJrhslkcemtq3ZaW2qzTa9amlpp6IS
9PfYBVYz4bMN7//hiinhUJRfcHKi+ydv5OOErnIGWZ0iFFj0zamwSl/eJztE8c/o
R8sNWOo5+kj7FhB2dNlWMcSfzndhoR8SqVopG+uoeWAOS2IsmQ7TkIemsfvRtw9e
qhNceVICC25zaPz3EjcJ6S20XMCCQs248xEeA6hh6u8txOTXdXqdPi2Gyu6Ddd3R
LgkNEm5KV1oxMuqEqZQLUKjYU+BRvCuf+gqFIilqyPqhFmE443V8DXdPIDyfpn7F
MuMrwbfopJSQKKtkoFliOlOMNEbjJxjd6KspI9mPA8wh7UxPj3b2RrtjA2LIduOU
kvXcsvvYTmgXcRRaLNnwuCAWn8RMQG/mtHpe3/4fOjatIVWr9POO0RT9KlpngWqv
LfXuucPuq06NrgSLBzfgoQ55Bf4GP/qj4jesyvtNq4iLQ5qcliA37G0QahGjnJ8T
RvrwlBqgOaXrEntdBlmTm7ngsx+rNpm6SXakC4sNS574UnVa2hAvp9n7ZTKzPXwn
60YfeCS9zc49uEtr33mPMTN5FYapi1AYki9CFxgKjxydzWTTJM2g6JHVwvKLMxTp
7kPzHwlmt18rstWEfqmaaRGAzk3ANGcPBsl3BjaJCrlLOAVYqyQ+Gbuc/1xuVwz5
z1yO3BgFc5xYBX2kCbaeGE0cbBWpC4qdO+Uh/iyBT8G2KJudPY7t+xArQCADEOiE
/FQx+GHORwqMXEmO2ZDyqRuPjL/ws/U9KRTMzmk/XqbZnFDwo5rXwLDbsClhT1Qk
yOZLR4/OM5cyGgey5Ywn0asPEy3IYJrgFRm7QD41SQHCRjpcgYgVDGv8JL60WAdG
TDphWF0GBd5ieiluVjb/uLC4Prf4T6PDDxnA1IUbTJPEW3yjv6BQTbEG3odJJc/4
KUS5cY/vfxKimClaDfxIWoGTPJCKEXRd+mVCzyLn/FhokDTKJK0wmP81V5O1oOZu
AOKYgK9oa4dKmCQO3LNEyYQ82NomA/ejMUSN6d0BqfWADV03yYfH+DHUo/OZSjR5
PjJYZCTMVJW1MlbiROuU0EZLft9ZdZ9/B3LLxC+jNtTEx+7Q5bSyR5k3HLc5+qAr
38Dw1HP+0lAGtwNFYaMV1GJyOCpbRIK+zq8ybsEo1ME6PPXC37uEt6YDqh72nfLa
pw7Pkog+EqUSJzcznvUyPk07QAac81EgIcewYrWViEppq8ZbU7WIzNdZqlXXQpVr
gswxZCu9slsnke6rtpIsw1UBxL5qR9vLX/1wkRVGwXeiMk39E2qb+8wkUYfTPA8W
NdvnqASma12CKLwF/qyK199bkeySkicWsVTfouOQe6zOBjW2VajFKpvb2OPXC38T
MQVyq9SDCw8OgnQQkXaPOOFfwytr4FzXKHsmKzqnsoci8JKM1ZmJX/LyMPtoNQh3
+J0nagPZ4M5BFpP61mSyQVwub1+g+7MA4FZyn3SBqCEqbTHeh+edkuVc61NBwFTk
QltbYHiULMnsPKconIl6dPojLalCe6U8WGw38rvIRG9pVTeXr/pJ9ZKMvHNG8T7q
CbVGKWrg7QVUgV0sm33x88COXYt7/YCql0hk+wReV5sLSfngu5dHnTxuIOb7h1sd
wnypD54gn8C0caJ9LUA5S3qvuXzNNRrpxRpTGKFAFeTUY/x/j0kk8sm3Kmng5wMc
+frH7sjnVOu0e/Q3HausH5tgYPGe4AfQa2lc4I1ey6gdwMr8TB/4p+mgYoXUvi5K
4Mx77+Bg48d09gJ5z4cgrBmZNz0lDCFo2neO4Lk4/mg6JBcG+7s2kaiVyjHAmBFL
/ek4tjOsLMnvlhFGRbFHx0nQyBQcLyA8aSmz4358eDL7UHqINosgKszzssoEt75w
wde622tA/NeOG5Rkqs+xxpiB8WXVch69Nc5Po/WIHtITTPMGzEx6h7e4zf0l4Voq
9By15qWCIcDi9yuF6juIZqk0fEQBLphSuF1dcz7+s0UInIBbOZXR+foXmjEG9LyQ
Y0XQB1zmy0CLwtLlnCHpG8YfLVEX0e97r/85VRopjeI51np8citd1Ne+jH0T3sXO
jg3R/pi3/dc+S3i8ICdvFChdyz2yxK66xlbKd8AqwZEtImVZQHwerrESbKf0CeFO
7CCwf6Sia6uaMh8Jpexig5KOZEGYhb4yqpTtRxKLoyvaJITLL1Pnta39x76cgjX7
Q+QBnFZ9j4sUPKFS4x3n78iWs08oC8ahZ+9gDQWkSUK0JV7lQV4knxRYQA+2CrZj
57viE9YkkPrt5YzXqkk4uZumlWXKUaCXV1JI1gYUjmYG/dpZlN3zugfwmrYybuMG
7gWTrYZfnrg+RUk6CIeW3itvDNit7sBO0dgDm8M36UjikAtBP2i+jmL6DXvEfMN9
OaY+r88r8E4smrbYa9K6zWwmPkPHaYB76YjFQocGvkN0IhBvuh2+OH0xfCOUoKJ+
6zLMNnDI0L3xcxIXzmAXaEO0sbeFyavl1UKVrHeiJ0V3c1jqmAxoRR2gSBN249n5
kUye8YHiT0Vhwl6dOjvyDeAyyXlCLZ+LH0YM+SNKX9v/MZSdXd6QLatuljGkSQSm
j9a2evxaRUPLeosNpUgmDfZFPbLokgNOy/s8L7W04CsKzz6Wsvln+XABw1xEN7pF
qGYoxTmhIVdirn869BDFRA==
`pragma protect end_protected
