-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
CD83zaBuH7EibhwBfGf+za811s8FZCImM8DPfYA+PWW3mgq2/K/4epa2jgBJlxfr
f31ZJE9aaisiYAJdJsfRYaN83GU4oxyv+h1VBGWpAQV252sy4lggyCIwqqjFUzHq
Aem1zcjYXNQEJ3106/MX7dO46mPAyCjstVm3dQnpVMw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 7456)

`protect DATA_BLOCK
dX9YIoCwMzeqIcD4Z7RRPGFXwtsQTtvbpma8hfOrk58hgyRExavPGiCGYuAzDUS1
ItPuoV3vmRRbd1xks5YtRovDiulK5OedojzYQG6QwEE2QOnCnM1sa7BTNh/RJLKI
BDPETz5kwDaxYEANBr3/xtyriVBf0uirjd4JP/0CznbmVtFFqI35MNrDgkquxD6X
ksqz8xlCq5gOz07ztbS8jA0qy07L9ybVHKFR1I2YbOQKtFJfxfpA9LUYngCH8L7k
amQFWzCo32WUTpE4Sn1pw+unOJHKlBZ7HHayoucHtww4eoZ++YLy9uOk9gkOoCj0
YMrP4aprbTDlWz7S6eP2zmeVve0H/bsr1Uh1XpvqXHEymlBjPPLwE1iAmTPx+0YI
CcRQX2D2Keg78rjXtfPoyBjK3Xh9aoxYX/dZl9p3DEWmn7QN0Oj9fjymXGPxOG4N
UTeU4Lfltf3MLXFqacI5T6gF7jTONk0JSl61T+Ka8bxA5Zv+osRAUvI5Bqksrt/l
kD/qSzbUOTToGpIRb3O64/mKcAxQKgZqKHqYfQ2ZrO2qYlC9Z/fgSd44ma7oqTT3
ruTaqwY1x38tPv14xfiei5gkNM7M3MRlWyRMUbb/MacIqnp1XpTMq0zXoKm5eglC
StFVDM8MrIlbX3nI4Zm5wyuecG/0UkMXFCerVBi2BQs8j7KQslWcn/OkwPNDoBGp
IBPczyEnZ3uwbcQQ9WncGx0s5OL6Mrc5f1isfGMpfd8kMIGAaZM1C+gIA/uIZug9
s1l+OErgRVWQEZEFZ9bC7yBIGEVdORPOX/KKSg2amQDqd8IuB2kbq5MpWWDEOxzv
7VVp99G1iKNiMxJFwzbcUnGoyn2noMKemq6KFMMF4SfbO+oIP2nxvojRBThD0mpK
7Bh/LzNbXoNoQhgqHwpoiOR+/aL8Un1uB6VyhLZwKm2/HHGX5Xk+atEtfm+CFgFN
5Xvriwf2MP81Av/Xt8oqk5gOFLOguE/Tlg6nGCwPDwOxGaHtbj12bx6BhCOziOC/
RdpCx1BsLp8X8bF7XnT12Ijl/MgIOwHAkXAU+Sg+E17L9YblUgwsL93RA+X4ykkZ
yUQAwuKypO6EmBYZwuVJ9C8JRH9BRt71OPgiVEy7YTuHkkt02odtqLlzN0R9gIf5
cp0cB/BqpTdAS85zqBKDq72a96fpq4dABi73sD1DnF1GpBtk975xiS6LyN3ByGZv
kBjeH+MF9VjA7eKio6hVFzMMVtHRJVUTY+YyarhbQ3wvlh9/+uV0dPBguocBt0t0
Go4lhGSb65yQAqRYe9ObeShxN6hepcChegYIGehSEK6X/VEgogh7PN7B43sObDCv
2DpUDjsgnMAnNi4nciXljaqUbH3fPtytIPBv/7zWWaEjaDSibEP/Wg0N/9xg3J17
wZpbHppjBt8iUL+aYYJqkdranf+5A56vKIH3ju6xwas71CO53z8SG7+h5PA4jyUD
xnzsEOsp8B4dSHcxA/sTw3rJgj/rEC4c30JxFIbaPEb5mpwZRpUKEEW8lcunWmlC
kv5tte0yx4vNQYmJCVsT5LR6XzRM3rZxiJ3dR6eQsNcoYh1QuiMGdrsjYLq+2GVA
IlPVGI6JPtmAOhLylmYzE/NcdyMjPrSw4D5sLn/W835XuwTThl8g/NGUeg/ei7NU
fUKY954H4XG4I/A7b/1TkuelgYUxKPhDqPY3FLpqLNlelPw4fC0xC5NUTuYy/oKJ
4t1K2jEIQkEBcbF437JhClbo/qzErC79zIzLN+ru65rI4EAwZGvDYlfQ1e38rHMm
ICuqm4nNsHsIb/OKCFgH0YryQ2GYHaqRIZm47Sjs5z2NCa6xdJcNf3XyWH99IMSD
CVtcQwcpDMWU+BMdIHUs8X2XI/o70zrsMjQwd++iRE9u1l/0OuvuTPKsSUskhRDc
3OtKDb/iquzga40k6g/MwCycls6rxNIbMoF7pkRVW0xaR38x2LFGXeP6hlZrt8AO
gMVdc36SaZGY0KqErX+02SQ/Y67Y+xr1UiErlN0ZkVMi7XpjLkSILEhAkKUl0mUn
Mh7i+9y4xV4Dyd6jGpdXpzSAW2lqn7lnzYrimYpHIFd/4sN0zshJwAU7ZMePl26o
6AbpJMHXSYiQ2YZ8HH6Qh6Vzi19ZRMvi6IaQbauZge/Zmtq4FRUhEQQIYOPrgzkw
3rUUUsRj5y+KWz9WNz6kmJS74MVRo1XToWq3+5NkSom273ptvKg0dr37N/Y8I/ii
eq+LDY124jiCwqHuGMzXHF44HyrJhPauEHZY7cZtRE8/G3jfigKjJn5y6eRMmf5Q
7DCRz8Rp7AGeRyn1coS6MOH3Nl2Kn2+ImhNGPqFZFCZbTFqayRs3c6x2iFMRr/jI
rP24YCG1JFeR6AtPg3pJ4IwiccSpRmmRpyIhjs0H/KtYUm4t2aA9VQlGVipV2bcN
ZTgn9fQTliV+Uz3+wxIfC+ZZFLI0Y0Mso2mcX+e0KRP6QRY0//heZ1cgzVOg+yPi
7/lKley1Sy0h6vcqzQjsgPWaLLGfDZZBfy3Hx8c5bfCd/8EaPZuKeLUOx4vzulGB
SMfC9byd6TWSDKP4QZtB1CXUS4QgmPHZfkEoacitAWjVYN0/eeHMkscqMczzaIh1
CAOXxiJXjstKV8gtOFuylIrNpfaRyQuQp7plOeoZlpfYm6++WcBV1nCmYrzAFx4H
tdCiAwDSOMVbcoCA1z8TWow4tV2gYK6czg3RTWLDZN+SbJvMNIEmLKLjPVGppMgV
ziyp7FQEz7NKzC13PhvLB5JBzTfVUhU0NW4EeRC7JM6OlH+aXMFf6jzfJVQfnPjK
+tdFk+5b0bAT5N5C7igG9U44r+Nrj/Us2Hh0ASVRTNe6izlKhlCappbJ+9Zparbq
oNBqKUg1QbN2phQxJbBySPEavjjweRIPzEx5wwJJ5GdkdjJs0F9UMi0k4f2rz9DL
aXq27JnByGQ8Wjz2k5KB/ENdz5p/IWr/gxgzRWNzqSuYCVU8pL9wSuzQi7I5NdPx
q3QUDmBaRNYyLwQyIJbzanM+woYAvPJDXBpvd07suwB7ye7ec46cAqo1Va7fP2kf
mImlLWxhKp7VKNV9SXCl69hmGBGmrYZ0gyLc7e5jOn47E1lI3xbaV4Qqm6gjw00E
1QHN1qcB69SugXWAgxK4tpwV6o1JOt1WcRyJEI4K7CIoNk08vwI2AaGekUsr6uhw
Z1MYB/avBcG+HX/jxhXXsc4AA8icVbxRUfUM8eXAvRrJIFFYGyoyud4F++vIvIMt
wFhkRFh2SZ6oL6GuHb45DqArpYDY2OgWeeehLLaYYln0y5qTAMxMrCv0mN8306t9
CuFJhPyzdYNI0NHxsJjzEUuwo8aUcxX+991knSku5rxP5o5n1AltNTfDU5xtoYTX
4Vlbl4Kvg6kjlNOrWJ56uAFKaP7qCe0b9iWhKe/EC4Lk2Z7R4zb+WfjGSAIJS0lL
PpBfFy+wCWgkUbtdAuf4MXATulu1ZtNTR13HTARmBijGmsPHy32oPFDQkZm319RD
a78XqD7rbHLqcv+ZnZVLcKdZ7OPI6SCGkJJ18fho9Yh4IjZpZV3KLkWIywscGzxk
bq5rO8x8bhtgwStK7crFmcYEeu6Ke2fTs9zApK7YtgoI7sJnV3R1GdXK5H4THY8H
WFYNyvRg3tEqyIEX/4bVcFUccCeqRFUXUT6gSXELONRfLk4Wnndm259WYc1iRVl5
Nr+FkbUWTWXKMVk/zC/qaxkcMhAG4m2dZ5P0asn9y4UXFA1wPqR7rxv7Ha988+7F
l76PxaJL3QwSDbK/Leapv267oG//zOujpHsg+UAVEuP0MivFYazRd0HnMELJ0cBq
aLo+nLMEwLiHeleKxXpHLUWSIlfkQ6T8AAmA/NVExoUTVPnAhfNqC/bEAOCr/acP
aMh+VNSgokpJ0Ctlt2WERXzpVReov1ciJ03KlEkgAkAmh5HQRhRsepyPOlWpHxsI
Xj272KriS5kZorvfzcvlMj8KgTgtn9lTnAsDg5R2EyfOOjwPgk2EUAy3mrl9VXL4
ryoZiZlOfKTlAXaWFrl2Sb6O7hs8vHpcA4hy21CTTf3qp1jXmwdozXeoilkOtguI
sZTBKTfKNteYaWpMB3oShA9WaiwRkMhBbSGNMuUfSOOoAsM+fYy672l2WJkRfHvJ
0lthPWHWUd8pzLOt/sA93xpn1VVRqMtIFAuGpCNsF5AMzLJteqHTTr48hQgEGT0m
l4ePqXDTOUPUQV7qLhgIvmJBOHN8nJ74cbADDmngKMD5ohabatOB0v91+HkJDaCU
UwpoJWl1ZI21bRxGrwLqJLPFNS1Gs0PIxPSLY/O64p2Ahfw4RNLqeeCjZZ+rT1o/
WFGdPT1dov6DaVKrbcVzf8p0/U1f4euilPUAfzmcl+GapUEJYUoUZX63Tum+3v5M
gtv2GFy3Ta0bcueKpncdZ8vrYTUNTcursNYe9l07jIDRouCiFYv9KD+6IEy0EEuq
umnoA8vk/zXLYqd7ZGtTH1LhtbLYxWYTSjnaeCHywM4fxi0TvsQ8T4A72rN/a5Ox
lufk459ALxFFM/4vnGxQnz7H7DYVLfMgAzS1Fl7OMLHUbYwen2k5kqAsAcfMGzMi
Q8NyYTXvdGjUgSTSX5IYJBJUMvge5DpNcAQAK7CZUGuxbouS1d+3Oty0nnqVBfrg
ZgU61IbOa2PFNBM1GglW0q4ls4QxGLEymURrhZUhagpjHtLwYJ1nWayktNMXG0oV
H+KURf/CCBPjJhziIcHWQQULgBYuyNQpm7hzeCQxRk6X7ONz0yLYk58k8F2uyRm0
5V3MM+9IeTFtClFiyAQZS3qw88gien30bO7GE7dHyhshy43E4UZu0EqmT2xY/gkm
dGpVtLWg2lxAEBiOUdvtPn7qbpiNWCK6JF/pC5g6FmKPD613NnCEIIXPNWwqRB1x
7hwk/T4lvFPuHWgbQbCv6C/5IIp+oblXNBeyLXWBybi0lW0EEBrkkk+9y5VOrGDp
lBq0VQDWWHf74r7cmyKBa5VNmbQ7dc4dZhlg8DQ6m+wkBh2J9xjQIS6Ug/SfD6RR
LM+8QXxuhghlzp5zClFj7sAefVcV+3Y0/aDCTfr6dsYNOhTFmtQNmJgPUj+vz4Dl
EIHwDCRN4iQN39ZOVOErHuoOHkfA0tEcM50SqZ1rcGe/en11/XT+TopvKq+de15N
WP1w1sQey5SLRE4K+mKEqeqUz4k4TRjXFTWW7A3YHEcWcFL/nkvLvXcrqFYc1anl
Sh1VP4Cue/R542G5wuLwMGmo/gYPp23AFEpEDS5v3gYVLr9XyfEIQ4HEP3m1CFyV
WnmyjWzxrodO5U8PAysZExE/malsBAEcZApT+q4+XGcBPHl99yV6+b7Lv7VI2Ues
V0G2HvcGlxI2LRzg5kn1HxGVoghoLiM4TA7/YQnjkzNI16wXdcYju5MymdP7brRT
pny2TA87zGtvEuPcqlGZtzaIA8J4cNxBnE9Wrosfo0D1OfAwB98mtfEEKn5TUYQK
IVD41ynpNbCAz62G7YlVXdZ5UokmkP4CTd1ALHhXZZATj4WzPZ9mvReBfO4e9jdS
st21/JRVOKZpwVn1GNjT5duoHdWEnjYHZDvRaeeUm0UM2/3l7EMZvvUXY2ID+joX
AdtRIovIAlDk7cyEUINiREOMk6DPCxknjcbH8kfliECj0trvhc4YH7sdjxO8e1Ux
Uj6TbM1M8IWN0U8ltO2SA9KnHrTnddiIX6/Y3ZmEx91pgVqa58HqvCt5Ovgn5k4D
ZYivEp2nxja23Acxg0NRlqzPQX4RiLAHeGWbblU9nbLSp1mKB5ah1cI9e3nL3xeA
7DgQb3nKw2mXKmBLA7ZBEILUWss8QHeIr+/RPuehu/+/w1wUFmZwy429CgCpUa9/
oiFY4rH240GC8hONgt4Z+bYwIemASQ+qkVPrPWm3N7J6GkLwo+8m9O3ubPJpibiI
iRLK0JCGtgC1gF4SggrYs0Kxt/Q4WXeTwtVBNMj0anUsFPZBSo587xNjflOqO8v6
PzZvTBIGRaEmfA/NOTIEiTpj44EpI+KxutZaBAEewIPrYjaqnisVsoBCDtYFiv1H
4ExQ5lJKP7OJ8gWcEwfi5Lzy4sBVmMbEFRUEDduErhJ3FnhQnOmFfZW2zooo3oaR
b7WeS/sP9jT92V3EO5M64OiJJyY+dGbybGzv3RuAbiOWrSq4lAgC2inBb63Zs9cE
G5MkCsoaKURNs2FJIspIZiz3IXJZwyPhWZkdO2i5+zBIP0858LhKgMzJUj5B+uIo
o04TFYDqZFaCsKFLb/6+90PUQNaQI8PSJwxhbFlKjvLHBY39KAOxIiTWJjqI/PDI
umMPpqvrlqTUp5uRTj60hC4uVpRaCoNnTvK1zRpS9J49OyRtERi8vwygzmwsINo+
fcueFJFsVP6DmkMmQVEj3Dg/sfFe4jDo6mXnVH+ehnUYQw5/fnSRA3H60mH8a30v
XmPl/BfnppTCdydAvoaytoAhKxdvuENMVqeQT7FAqvhzTKas2TwPcGoGE5GQCnmr
9ptVUMIlLfsyvBimQ6KmzVoVd1+jSEOeU3uOWxGMPTTCZCwZSzgtIQfiRSX9EM8R
6OfAo4cP1CijNTUKvyltWRDRAzY5D6iWI74aLXxlfDIAimzbyAe2ric3iLZLt11T
OD48bVFxNklGsBYEDhAz5qbxVGZlYWVxa7ZUoW8HfEo1NfA0GLeQJc57ZNOPxVwR
gJV/AKEBjLdoyc2T2T46aPGyvfu4qjH65yO2PxgDo9LT1QVc5u2jKZQoEkVt+CEd
AeeRFL6QF64nQ5Ax0eBm+yHawRe3yIZ0WgkT0xIcMQqWP39eZhIcfxuPV6ckmpcZ
gcp2ci2yiS5TW1zJqaSeTiEUGeilDeiHhGyEDQuy8ZgEzADb8URZiJbUU+cNpSJK
rPTfAG/0y3hJSnzV+stBGvdAww8fJF4OPaT8ceH2bYUXaexuIWsgHJM3SzPbsqzc
tLfAblGo32rrKhYOlXqe4PSwo1NQsUzaZyFdKBttnLid0G7jpU8ntdnoIQVY4dYP
ehI6TAviGIQAJOrnjzJRZgu/bIsHqDmxvS7HF1YRNOcZDXZ4z2dDihvUiUAZH98f
NU+qnm0MGBOnPWicq4R1VN9sD7gYb+FptLE3InurGMVclPo3opVK1OjkcuSd54v3
qeWyUlj4yZJyMtF4B+Vl9onKUNb63eo3t6RaWhICb45x6tk79WmkkFWJ0WvSmXWk
Lva5K1g5nC1Fdwolka3m+k0DMJlHxnmar8pu3KSjiJqrRSEWkBiPACbquBjBgRY5
ib5qOwp2UUh43UU44g9qywlLYobyAbRLeTJGOnT6JmgKndHrJtlu0I7cKG4qcpKl
goKuxMDOW5blbq08ttq3e+2cy5/bEIiWTn9MuulxKogIJ4m68w/NsX+FF2RMJazJ
3zaxIKiSDP0vEk9HcpZLTN0EWju7NjKadUVpe+/Qbjh9YDkwS5Mu/bcno9k3RE41
aYElY1N4zm1QAIOU+f39bSCwbBdHMp8l++fMIIMvHZStDTP3o2SBiDAUGh4/e+sh
lGK7n+3ccyiCbGf3K7OSRWKvf0D24oKvy/FRPewFOA5XTdqdkaB5p5sLE5DJjt8b
mGQFC2J5/t5rN3k04xFX7SlefPqvXr90ku8Q6+tfgPTkuG1JKbpM/vxbHnuHcek8
+r/7mqd85tnZ+Cg6OcE9PBKQR53xHN+7+Fh5iZPZjVJz2YN0aLEfepPrZ82bpxPg
z7nbrKvpAz3BK1qI+KbMc/069GP5bmUTfeLzpCOgbu8/Da2Px7EEs2Ji/TFlrtrY
TvW1DlVZzBlvoJ8PQZA7Y0+6HKvScyZYJCM/ym1k7rmEv0RVGtC5hUUNrdMI72LS
w3vpQVZsej/28JpgM+idGmWfe3I13xElq02sDDxWHdjMTrQV101Y6xo9rByfvQWu
Bm+GyUEaFdKLL5itkyEHX5WvvbXmqBj776TgJdGfFg0yKDxRJKUeHLMHW2M9uNkQ
mZ3zmiHjQoxg9HdygGBt6mcrK4woPd7QqCePNFCrhWfE00N/SpLIrELwO4pDJFw5
0/pdNDDZmqEwESBPvmvEJKmy40zJHg3X7oRIuAaNGJPJi32+FpiuxGhp1hp99lF5
J+zfBMcFfeINw9eXbEP9CTgot8HKJ2T38R5kJNwIju7EYzPKtGH9D5tDNFyUui+f
qJBz9/qApZsGv7xH4zJTjw0CRwOAdnGW3W0hk2y4LD3jZJuif21B/tv5KV+IZXOh
zlkXYbvfyvg5Y2AQpYkBSJDecCbe9Ck2yidnF3Lays1lXzU9Q9EuqU1DcUYj1UJ0
ACcSwOGqJOlFM1a+E+a2O7D1plhQP+Rzy4PXeA/TYgPnzKZ72jdiwXQPRMlZOP6/
6iGTjgLb4cG+9chyjRlrlZ73T5Rmcjz9FUCWmpcJTopmG1ISDRUKJrbcARWp65M7
vIM2IxidLDJl+GDmrszfZWLc+iGWnTDfqlfR+XNsgwDNYjDo3R5pD66pQLcg4YGp
IRfdBZjVrSLlCgaHWNIuJm1GYThNAQ0nQuza3mlITLzkfA/P0zQ9l5kojVVNYRk0
2hiw5niOZPCAHP8jSh/XalFzL0wWyNujq9YLdfgw/DwZAex5J+TzeoN/HiGP+TvV
7gEV6BbPNV7JWND9r3Yvr6N6wzSZRDsmrU9+RmH/3pExLxTS3Ff1dLQMEWS4BErN
zXmmAX9o+kIPtrOsDUDujnV/TH2jkaM4N4oko1uYl3UoViR8eVSvbdFfMgMXCxin
SLY8Bd8KC16CNSNFkVFJcgVj1MvahDWb7bzuND4BgPhhnW3HhkLkDxD+/rvO/TvM
HthCkPXoozNpt9BFv7NWxSauJ0iIQKWXneDVuJj+ZSdb9yzn7N6P6kYtrL74UokA
FpSAFV8xY9mF5E/ltb3sfjHEi9ScPopx9bwk8Bn6QDmlkaHNAT+UPmx8S15wKWHj
eBBN+ypNCXtdr+9WzxMJ2qjz14nleHVeu5e/hclnvqHdYlrIs+V+y2sptoMhVttd
Vo2Ikqa6Gw8NrKkkFIUkam8VySr8zXnMgQAc+ZfKauHu6NMHfAelKSph9Zckv/zc
8+Bi23XTmJjxWNihBy9L+D5ybDBbimsBba+nKvK+K8ZfhFiEkBSXMUD2krhgW5XA
8x2+Ol8Ok6pkFw/vo0WEMGc3yIml049JyGXhMfFkBf5B8hXbpl8BFe1ipbbPAB7F
EvoajtMkmtPsk2lSvFZsyyhWx+vuvuyURtkbvVS8uWd+giQ8cikI2ZHIN8iI/g5l
9K3vLBP7XrczTKc2n9zvpmxEUNVYVq2mrPLPHZHNz3OQw0dORu5R5gofmb8dasM4
+zGQiQMOGHaFoTBT6F7YVdGHCizhYPM0UlzDDt37Aix3+jXILVB7RNjuVB77BZqU
mgePLkasb4NolHR0YumpT9/YNTKy5Eni4qIsR0o9xGR+Q1pwq0aLA2ZjnRjiOhn5
FJLqz7ZlFydgpS7Bkru0jkkhPuoYZZ4MRfpaNOiWspUm39/jKlD5kOkMC4xIdJiU
1xe4HuGVA3HP41Kn1kWVCDlaQR7TUZrawes1HtXuVdxAsKjoSWZOF5gYM8jwYJB0
lkRy0/u/k6UHXZAf0PNVDubYJ6DZqf3ZkjwH0txlZinraC+ioyzHPJkBUUw2qxBN
9gMDOJqujdx4T2wkBUn+gZoNaYTEEBElTUscaFdfzzqwdvHIZPmszoG2U+8P01d7
5qLoXud7Bov0alGTWPCy0Ef9IIt+dQqBQCWyB9NobozRiplJ0BiQ8++aJSVeAlJq
0Wei36urmPWIzDF8h7U9G64MZH/ahx7TzjS9I5x58D9fgqYa/cS8YgGBwkqPnbof
Oc+V91/6YI0CiMiSrVNviCeeLXIwrz0JIOxmY3XRUj4ffvTtpymJEFw19qvmflWS
IXHc8CYLpZV+wtS9ehruA1fZ18sZisjMV7y5PEkhg+bByeo3QTbN0V0V5clKNAQb
`protect END_PROTECTED