// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Sun Sep 22 20:49:28 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VM5HJEOPB0i3TXEdxXzFr5VTq6EcIPDZujJWGAK1aCbLXG/2y2dKNkizcGATmDyZ
7xVxbMM7FIVsFPXg6Yur/Gvk24I9TAP00cL050yHcDS9+YK4zNRvO9KwBbuFO1/e
MJpiYf9rerXynDOxPHSfVSLEpKM3H9RxkhcAeieis5I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23792)
+U2QD+JATy6QdI4mtJ/iz76w6lasir6jC+5NVwjKEtLe42TdUIgNzYYayXVybjFE
TMzYgtW4/hp85eucgMPsVz4NdBM41nmU6v7XDrF8AuZL+CQjBGJJ0xj+kG+meOm2
gz9geJOXT036cTlMuFF4eQtY9BAbk/rbrvJnU7t9LnotWHB7dWk6Jy736UltMmO0
ILt7eyDnbEcA6yGq/lX9em1faM1PuVz9zm16c8+gi3KmzyljSn6rXC2AcGO+Mb61
Bw/X5hhVD/yKGwaqA68N+FUfLZsZJh24eL1nDkeKCX6PvbBXVGsv0fiFdxh6tz42
BILs9z/uBTXA94Sz2EgY+dkPALd0gtGKuwZptavmckanovX5OMFVJ2WvSJYworcE
988v3w69S3IY3r0hVDPa9HHDaoUBWVl1jwu+PvrzVJtsrufRHxnYzhOVCehHhl/k
AOBpRilgHdZ2VHKfrWKPbkiVDQeXwVoaJVnH+I/mzYrsgnYTJ27S2f4M0DGEpNHd
SgqyxA8+2uq5tvEx8lvoFMCiE5RCk820BjKP2WCOiTRbjQFb9ysvZoj0s4ppqwvn
1KIcfho1KiGwf1eM5IUjSHFqD3U3bjdhWwmp/mWpgMuTPUpHsLuYBF1XtKGjYFCa
EBFkRFDjt7TT572+XU9S1s4ukbu2o8EjSqXf0k/c+uko8jcLjfDa+JlwSym+dymq
NvV6gzJ4zqiEqQsMhikFAEq9BFzi7f7bpVbjs2MaOjqV1d+r/xMcvDdjyEZUnTGL
iQu/EkXLqLj3JZ/fj+zrMcC0jDnligHg94PVc9udBtn5zj7KG4PMm8VSCzoHi51b
mw5TIeV963b5kOA6f4iDZCecNThzmz3HbOmzQs0YnFV1rLbFHNUnQK+++IafR9jk
x9QGf6n6mJFwwO/sBPTQ5Mx1e3cKz96Hw3cXMkajGEfR+NHBzgDvkQY5aVttcvHa
qcP4uMnDxuOT5EqOp6AVEs+6QxnnbnzxslGBPQfWd/MwYxU0bem2Y5DEQMtVgMZf
dca2G8pkk13DxQI18+UA80CcEjpKemabKAGRw3kDeZKkD1QJeHHfTSpJPSsi77Jp
vKTsIqbOSDWgS70KYlHKLPbszososZZXboPaOOIZAnwDcC07qQOiLQUmFQoX/DnV
dKXm75D5JbUlftYJBiASWiYv+2LVPiOVokycUaix4XGIlLObiq3HCe/eeBuHcV/C
0J9hdNrk0CPvDahLyRTd0t5cfSFsgyNs31Aep1lPgQ3aiL8mDhnJkaVkznQiO7cx
doIXw3mDeT4dg/RdwQynmQcbIesMzeO9zc9gpsi56zx0ZRUuOn9ZLcoGnP/T1kym
Gl1H2AS/+eubw3OHKgnUQQLcgFhxpYH1NaYOTXVx8iKRsToJD/sSS071VToDd+Aa
5OeBFBX2heKQb7YvO6+WZ5F2gEbzHK8mAmtWDiIvL/vRbal8q/k7HdBRicpI9OeO
EtotqufQ90MMnFBYM6NYBKM6qCjBlGkSt0iDrpLAviE7mnj/0wgCbhbkdRYQde1s
QUPC2o/iz/7CJm0wYqZFJYsuVN5/eE0xbWEXZjjHrDZmod9fd7zfSjQb8f8Yps3r
VQRql0VKpFA267JncmeLJDZK6JnLlCcF4xhfngO/Kc4z2KX5i25G9OBNVotbMMs+
5B8Zdd2jAoy7vj/lduZrgpqSlkCGg3yoN5scBlnZZLkd/VACQa5peqnTjKXFE1sE
8CLFwD0upO/zJQvfsWQWS9YW6qmni8++y5IvkENtFPIcboVSXoyzHsBN1oeWWknx
k88SdRMaUwViaU+JYUc6UY44gDrD6FQT9PGwx+NY4p/J3cczIXEU25yeVoaZz8QI
Xol6oa7l3f6BMO5ZjDJrUPXNPqpK4eRn68nzmRYafbAuqOX6wTfpuW3LUQDyadPZ
Zz9jBLOCG3rzYuT7gozOk9DAJndMeaaAFcOWbO4PM35rRMRd35RH26kZ+yB42Zh4
8d99Nk0HqbMsKmQELfamN+MZgrdgm6B5Abx/VM5k4p8V+7rUVK6F4o/xFqtBvtyi
XdbsTPEFbb+PK9KNeXUwRH3YDnY3VOOOimJHZPlzp/fgLnfPvIR3Nm0zgV3XgsB7
eEeIWVt5Onz1ywWKgyf+GTQm1RWrWATywUS3djz7/bH5MyF5RlWEjbMYH8b95fIi
MP9gBpDFxA/HwEVyxBPDKhUxAeN/UNCB42AzALiRgPXHdee4Pc0RItch/tIZSzzs
1o+VLRN9pY6aHdljI4CDY+WQwJLeCjwFVMf3ZH5VG+b2x4J91/0wAUpROk8mcItX
g9y434NsRpaAN2/OjXU8N5TxBnLBGBk6nJ6qThdj6duzTRfJ+6U2w+oHbFp7XmV8
aOe1g3tACsu5PKq7qSiz2Xyz5lcEI3GEJVVurgbYVk3F2OUgVT3APEGIQiZPbtkl
EOiI+h6F7Eb0baMb+/jc+3md8K5XFfJzWlhujBnavHel7DkbMpw2aem7zMogeJ4h
KGKFlOFe/VnQDUkKjvNn6IkQwn8xiKJRG7fUPUi1b6R0YImv8YwX2E3FmDFvm2dX
E14H/u1iVbid9vBuEwBf3RxJOt9vW1hW4nX/zmoUNy8+h0OHnZUcOqJGw0ToVrTf
O/K8oIybB5W/UNSImza9ChjsjpWO/1j9CPFp5CpQDzitoHBRlKkVutRLZ2Dr8Cb4
HP+y/L1TTiVPr3Wt2oTB3H2Nn75YZtmRw5IdAD1KqbmSwiiwAe4+5ujncR7/CCHZ
kJNNSfOxM7FCechLBxknwBN37GqsRjpg9dxaF0WLYXc6ov3jBAKuXf3YDYzrIgyW
EjsSzLZe1Ao6BgWfahF5gKP1TgFgrqfdLVusiHetvcjtl83EZspVY9GUOaoHbYp6
GOE86RJLFsEUX0GSbKPoYKVL6AFQwIFTL8SgiqyNiHJ8vQTiCbrY8LHQTOGD54dt
suRfaZkM0iH0u7zums5WaRRKzDiUL3FVj6e/4P2v9Rbow0+SyEMvV3wVembJQ+Ek
1W2doWToQr141+kTeOcwO56XhHeZwicg6KhPNoHMeg0kToQpBqLfQx08FlL6ibO5
PvaxZquuFXE6K8m3OXqGT1Bu5opXVmn6ZOcUVYANkwFWaGqIuYLhrlWFxKSoIxv3
SJU4bRSVBrSNag3ocd3z414GfDyYFrLVGy9WEHSfAJZ/TWpFcgU8sO/JmguzpZHo
g1y1z6HgJM0DPHfJcVoMFoNJEZRaJx/+xgPEKETTD4pt9zF/FF5vvb+Ywxn0r6vs
6yX44CL2wbeB6g+jynWXIxHaSc3s1OZzRyeaN6TunOMyNnAvoCMsu8C8bnd9H6Mp
SEOSjR9v5q0z6oMl5LH3IZhf/OgF3dehUA1pRwOXlmUbuXJAxJdwLAgle9+2d7P4
d19OXL/FxdZiC72U2A35H0jqgH8g5iz5/sKClAlr/72ETZVdR0oz/hO5S3cptrQv
PKAy+xHvFO17igO8qaA6J7trtDrDzhNc3tg53kE4k0KmgudOFjnVOawi8snVcmkY
kbJ5SENMbMHFGhQGENahR95UQw/FiduemEbucPLmeb68zrv6KSL/QACoDKOOv9nS
54zEjL5frBvxmFTo00lLbMUOmsByKnqlcf0WdGXCvr+dVYGq5JwflcLHjRwc1rem
M1a+XlviDkw/2f1kFXmQvMPhSnHrmQQaBxlxBWieNLAqhLfo1a6TTwMjz+Yi2iwW
VtC0UjRfjKmm/RgTrAAtI8sorTEEM5/gpBYM0m4p3r/4vOzLanPF5On3PWMuPyOk
sLzmCnj+jNjeOjELxX2hQpLvoqrBIkbjlHZZjipIRrpCjNnNu0jzvfQmVKLQ3oh8
F3EzFW4wCCQonicMWMTveg8C4EpbZktoBQFzzesVrbGOSZmJDfiPV0GAUWt0Njqo
j2Mw0qSZYRH6VVx9fXjdbTfCvcEB5ns+ACYBLQGGgCTXcRgW9O3Ex09qHA/WY62j
ZOItJ4olwSKJMJKFuuOWkLtBsooGoGUFpSsIYjwTTjPj9by5BtI+QjpBV34oqAvo
KsTmremqy3rOEop4f46mxrPUKixc5depVIjhlkKkoI9wmrbIYbtYDou5tgR9dGgD
dyv7OeaUg1NoXqOmZ10yf7XYXN5bNj6snwM9MRASU0SzWg+FKl6GTIsnVhX+VeZf
FhrVKhyK8IE7OAfHjQE1CNY5NGU1X7Bb4BxuhB5CUm5wqzW2ubB8cXM01mNmqL1o
+g3Y01sAOgNBJpXgVXoAPEcIrJjE9aLqOh3PfuvEtQdbBC0dEBWupuIq1bXOgxLr
78awXwazCDlNhiovZJNTgJZ3AGCrTTgpPOxIXiCtV/sON+p6pvta2+YKTH/Bhfyk
ZrxIhsvjgsEmIQ6PMREiGclrkhknEK59XWEsPhRwp5bPjcOKo/DTif7/7zia1alc
CeJK6gWbwrWSiJba3NN3CRvfRLxllIsMJBBvSoKWl1KWjSeaH/RimdnkI5g4Mlvk
BmTh6xMG+AX01DJcj2znhRmD84sslssuXF3P8hP3luylcYj8KNjDtTPsmeOZuVMV
v6cLUi5fvfiQTWVxvljAyBnIhKj3kbGA6gP/cP0y1+2pllztiyMwxFfSq/Gnp2lN
rxu3Sor5YrCQ3I5GaFXia/SqcT2zlMda6Mv+wO0JMWhzsqhOR47ph+u8CYaUt87R
PvPkGAv5rvOCYVzzjZQFScwrQetypJtosPcIu/3g9AFMuXtqyg5e1a2io57inr0c
TIbM/Den92Rj35+CRU3nKxr2FSNqX9etl3dJCOm3o9+iyuo3ApogShGIEqLiM225
+UDQIu6qsQHdLysPhg8TgcfLHvJ4eAWBX3Qi2V9EWR/Lq3ptb5NlVDspylCJ9SDU
VcGrEhZkiikXjm26o8iuFwkLiVNKHp4RR2v/dk30LFHX/3/BR/qgUi5Cb1ONgjph
NVL35A5AE7KJXeDLwULHvY6zMe2b+zGF9jX8/LgvWeT4911CdeEjG8hpJ33Z2m2h
0UDr+ZxMZZpWcdxYy1z/FUIUASpmR4fztps8jumy/DMgGbskVhRZPW2oyXSlh41P
NJZt8Aupp+osmnVX5UxE5s4WihFknKc2+yGi2rFHcJjg3lL05/X6Bb4sWYk4rwE2
+brzj5xXipG1ClhbDwER4S8SbmdcH22MWoM6m8UMVERmM2MyEeBNR/gZIC8Pm2kC
lWj+3kIrT4m7Er5QYNnvF2jc6ye2vdRoOyfJHS9z/UKexl5kj+JBxuybOb3jYGtw
fUBxW0tls7C/JDNDBNICvyM5smP1RBNp808HjnxQt4HnjNR8IAqOFh1Htdi09Ao8
a1IEUqvun1bEOsRdOddpmJaSqy3ylOz9FNtjqgLoVroF1pR1XOvbWK376Hq9pbEM
T7aQ3qUojecnzCSEkLAURuCYF4bZzS6I+8gxxP4ahM4ZUJw3usX+APVJKmALoWWx
Lxn2rcxVfa62ycYB7sLf6kunLO3jJn2Yjgl3nYZVgDB1FZ9uzs5VcCSegjFkN9GG
PwEwHzoE4+OLegNgNw/tZoDHnPZr9f9HjNz1EeF8fD/c0N2RVCdv+oQR7kK/xZDd
Xat+yCVv+334Ig7N6CYjf5B7EmdNNmjo/eqjyS+kejJQlzPR156joDuQqhEE3rj+
o81PQ7RfxWyPLe5hMOfxeNqtYcyFU8pCqjldohv9Xx/l5ODzytHYqdRJiJnI3Mkh
7qtRJHtOjhSZ3d0/Y8G/ISI/976jgfe+X9GPs3SY1yyjRCzV3/ogszF+a3WCE/oG
V/CLfGaRI1/ePivTd9TB8j7FBcqioUvrKIYtbkZWzcr7jrWJcCJQ2sorJW8UFY46
hQk1gEQNBmQS2S0FXrdjs2WU4kagXbRfTLHjM2YQwy3/5xK39dtkH3BmTEbzQcJJ
kErgFs66WMO8BBGKxKkR/JnSInBBZqyeuHwJxHnUw8/VZMr6BcVllpu+ywoWiFvH
sqLmNXVBzjs8rAYPZqTAjJFi6RjlOtHLcS7Zb+RshMxokAscPohrDhpYz07qZf5Z
2OQasZOzaSYduT4HMxcZa3MAo3kKTd+zNAsCVnbR+gC1dJWrcW7RM4+PR4a2xxjr
vDmAjRfii2IOcAfMrhxupfmjQL3PnH/HyJ9WepTzdj7634WoKYnxilXaILqhgYKP
WcZffbaa/Bk37mZh3YpOLjR1bDU7Lgkk6JGME1+BeOiGVnpDPSdKsfP1gVDif18l
cii9e6KnYeiw3DmHFWgmTq/CKM5hx0f9n88cWzqMm/NatYgJCPvpTYhnay+jGTKj
6F6cdXasi70wIIyl3hy38fwxuAV4C1Ep0Tz30T+SXzmupOimqn1QCQIjZEalywiR
Hdrl3QqTNbkfNacOX5U+T6M7OUZv4/unT/DoU94o9BVDqDVbqk719LqGJWzk4EsL
rd2Spm4K7l0y2ExJUO2/yaN3FEEzpHq8IdafqljBnR+2Yji1cyP42aKVOxVOBP/z
kmi0ZZCzfHrBxHtyff8zZxr127uLKNT8TEB7wFkJQ5aAgn/qmsPIu5qaU/aY5qqC
F0E0MEaAU1frXyec9l54JdJZGfRnm3IoaZrekzvi4vaobWXjw/XemJvH5PaQQNLm
ESm9vLOUMoBkQ0TMwW4XDul9i4+lvsoGe0pQDYZCV3xQS38U+vQYHjHgRhn2QiAp
fXAQmiuQkupcvLUWf5WjVhzZOeGCnOaK53GDwQ0E92i2mF9t5Eol14SQ8cW0HML1
0YlTCNqJ2vJfqIZ9EVe85064Q1VqcICm+wJCTmgj6/2ZD4s8z/GU7lEspEvwLV5p
Rb/on+BRnbsaM3BuZZ3JedrTXbMkq0IpZX8z3x3FkrmLc5JQ65Vt0uNQfW1zDbuf
VHgpKCO4jtTQogWA3fJ03WI4okASIDqf3vFnLFqKsIIuoRkgZ+OZBHwzZw8b4Qii
WY8DbUdSvHcxsr9FhYbkfD1+0A5c7tQhw/VpizaUCKm1UeD42HRA4HJWHV4GTb3z
tk8dU1ZA2XuzFnDoQXDPrfzHuHPUw7yNjSdKyjOg7FfjB1QC1GBGJkxrW79zEpvc
BlXlrvPRSMm0cUbT3WbWqDLwCuREvJFaUlt6X0OIB7ZYXbJFd+9Py/gLyKd2yMuj
GVvP2tq4/oAlp1T080qEHOTqhf/DH2cxIgQ8UVk5/Ee6j7SkwCmJaDllkOWLIhVv
QDTcAIgUflqKC+x1aoI3mugrX0YlNk1UOmv23afWUZC7mnvhGS/ho2RkAEw61JiU
Lg3T2bECXs3VWFNmy2A1zxcMbeqd+AzN0sLOuX1sI567hev3IUf1n7JHNPVJDk4k
owIxTcEwj9UBE9b/ij8/fEaohsVc9rFrDjo6S50z0tdcA0vHrIDYITGYKUFyIlbT
maWfEPWDWzy4sFLARDHTq56NntGgziZEjlTK6QR3WDVGo/Tq/ylMlwUWrGac1dhj
Mw85yQ9+O4XhFJeAkQImqt38lKc0BhhD3zJqhoyOxACkDDk1k0KWECuYtfxlRNzi
e2WJKl0mZkwsK5ZkFbHNQcxG+9KArLFHdj/I78tDK4s2CeaYjVk/dvVtoONibShs
YA9CZZhKH6R6xU5smNGFIsursuKwSAf9bRuTmIyVI8aUPoBQt6/X0MqU5zLAzaX1
v0+u4E/DKNXO0lJH6cdMW3WHMjdMsI+vFIspI+ExKSqAx6PQQ8N7k1oTwT4Vq5mn
W+OEstmBIeUiwHU2YBvFj9z/urmEQnBfNmetb/cAKPhC4ZpB6I5IXmoqU1Mjyjnh
h76GpD3lNUWNvduUV9R2wOjesjz+/pki5aRMAJXXUMCBcV+tpkYMSModYqpNFste
C+mAIPqdV5XZpB1CBaxQux9iwX58HFFIxJfkOUXPAcaW2xlmTWSXyosXW1RLfc6R
+eQcoy9tA7bC2G/MmIkhyZ9NrfysZCV8h+O3xD/X4qK2cWY/4bl9zc1nMBu2gYsi
3wi3KQ/Wnwt7SqqIeOcFzRCgdsB2daqZoLU1SwPTskoQTDdZfaGsDa6X3DoArh9i
VCKpMb/qBvCgfZXF39Jk4GuIyw1FF3MSXbdSXSEkHV1YoSYuAp0eA4EVGaymQKtc
HlCuZqp78QQvOmblZ6CSVHcPGqQxiEgj4m51MeTEOCCpVGEkM+XfkyX3M/Eszxor
YtP8q0eQCKE6waSOjmmrg5y0aO/zD4EcuZavsgcbvDT7tjvVs/Mx4Xhlkhj1Amz+
Pl3g0WqC54ptrpXfjYgHaSQO+ZWm6sZYhSXyGLKri6FR6oOFKoqE5PwvSVxPypS7
b7rZCud87jlhF4m+mY1EZCXQhjmHnUwR/5+RKt3C+JMaXbEjuwVZnuKajVUfwo6q
bWpuPlGmwgvnL3k//W3vRZG8vtxCgdj07OwQ98a4BvA7LdWXCUPd2RKwqJd281Rs
j2T4GpOFP1aQeY7TKY0COWIloobzteArdtl/cRE+qe19vC794WUI2K9q4PXSAtro
3rrrLS2giT4NNTenOK+KSjnDxob7BoZ/GVTlTTvQhvUSx7jkp0jU6SGaqeV8Ywrg
EMQT06PJ+NFr+H6fhghaOyZSQwKoNEpM+1vTSpUV5DPOXgXNeN+tijM2/vSNkwoC
WCt6Fwfef/JKiochWoIdT7FeF0+yHkrEpLIq5IwTn9YdocR5lO0NNQhREzOpa4Mc
dOPh+lK/X618LHQiDs+QSKew4I3gLDMXZeD3F2ldWMA92a+8wwRmpGO92Vh9iawq
NQ2BKwKkxviCUZxTtYDy12Hui6LNtAKATn1Rqh4c6T3/8EyHikDX9PW8dHzXwStO
gg+fVg9elSKNUlwgk/zW++uOHNx01Q9DpPXP8SDbNlcVx7TzKFIE0IINhGAvxHgz
5eGhu+RxhZ+/JSkUPsc2X7LQbZHTSFCV27nr2IwJcoa94lcB7SAsLo/ixbwjupxL
Ygq9ZNf46j0dRxjEvc+luyh4kOXoDacMp+MDXHXTFnFTvJWBVi/bpmQOeK04BAAW
tBTORyA5rdqNnXwEKMzXkHxD8396awM/OaUxawrXKNBqAZzRrYonY7Athm2qY8NJ
clSElNpYRWSaqgjnOoBEa5YuUwAEvJHMlwP4FlEjn4MU2lhZtn4pIp/sHjVzne+F
lBMWZVb0Je1ny6H5ziGkyADYAMEAeSWN/IyJoDtTUNwXtp0XRheXKgIT+PLlpTs/
/OthcVDmNShirS6C3Dt2i3MKH+SNnXporPetzJ++Vtr2/Qv5tMXbziErG97e1wuJ
unJf92BeypBM3Cfi+rpegHLrumt2KtILSlGi5GGv6BFCxzviEpS/UF8t4rkh2toa
oAwkPSNET+s3iKB6Snqe7/6tOlv+s/WrwhmfifXbwqbhNzXAvifXzbTRyrklpWqd
W67vkhklrSm3TF+YXbpMfDswBu7xPdzlTrdBGHuadpmCwOjkXDdZ2CUvuDZK9jd0
MQ/eE6UVhDrkKxbU/AF2UiHJwYIwu6T0dGjWj/nsdFHYyM5jGcv65XhGdc14Vo3g
y0SVpxCwTn5R0K8e9Eiqu9vQoTQhT103p6bWrG81G1cZcGtylviv2Zls9Vq9elt/
z5Ck7317BgxRUXtOSV9A0PpWMYiL+ppENw8TC/7MlUtCsCCvMIx7nrYg12c8mkaT
D1y/WXvzZcX5FA1ihHmOYND9GnFs7x85tgGiqobmVoZ3RUJHLtWeNruKwl3FQJ+L
wTCvzmCovFFcsSNG3L2XBXmErhRmnad97+i80VemqRxyjvWk7F62WCv0ltgbNjRG
pTaGX709l1fsc+vr7hVxxdEbb0bG3/W9Bm6GiBwdWbqthIuBieiFndru3cW2mapj
r+GbYy0xnbRixY3CLZ4etM8laqjZ19AiVQQBl92szQ4kgrKW4epWuP5/Me5R2ODQ
3euqEPBuBaYaWkbhsGdkzoLEi9CTz87/wxd7xJ4nHdb2O/DpknMzSr1jnUGoasl9
ml+6D6kyesLiBlh+AQibMTBtwIyvOBplaLSJqrVwNILpS6f9xslFSCv2371dDHQz
TaKG/Mk1nuG/OS74F+XWsboWxVWiLLHKL85oW0iDRpGtM00DCWwjxNMPLhei91KU
7L1faH34uV/acGbAGzUFTa3FptQOtPdmgov0PV2ZTtDDteWp0p69ijtzOmcZdBIp
R/OZeX3dYtKnWKSdwAh1HEkciCkOqvXunYEEgJd6bjUOIBlCN2Psd7Ok4kGLSn+E
NwEj9hSlXDZB8T73J/5vm/a+ckjsBYgN7Me+cfQAP8X42/r200/R/fEv+8J6/ejs
5afz8mYFJ+2pY3CaFjMXTMJpi6SXvDu6xgaD+3VP0+j1KkaPcnvWR6ZZL7TVQbTc
zPGsJFKoGqzIjLMIWKhGPjosC0Eajh3Gwd4K1UZHMVbk1SOGUZCQU3G04kGLGEXu
KovG5AveH126GJVr15PsgMd96pnOs6Flr1Adw4gy5XxXGpGrnkFfwJ5hwUA3nzIE
jQ/n1kLXGkXanr5tDIbL7bNwiIi74DCwS0P2b4s+70waOwVgfc1dsG+gZCuXIqgA
5sR1F58RUjFi0dn9/F6IHnkKdOfnAmyrlo9rfDDRCYB+EsVEknuSlyCSt/GUdr3s
iE+0Jpeo87CDLXsF70+GWl4L+xviSvqP2CrFrmYosmeESpD8n6OOUbU1TrrQbN7+
LomFn8Ddk8wHYWSHY6vBJa1FarpwpeBTnJMiI4blJIiyPObDG7TzsG6V0B1yvwsn
TqzHGC2I4fVs+Lmsy5IPvzVw4Sn8mR9SkoTqBPXZcbai/g4FWDI8E+loMKJ72EvH
MYFshSfDQOXKoIi/TiyzJWcVJiCbAb6TVf+HfwMsbDc98deYpQMyV13GX14ES730
Ak7hr+ZnHxkpmSoNXGgN7Gq0U1gnBTgeRn9fcAYVbMAgsk/o6xYkVppNqBDapcQw
JOb5j2piWLGDF6ZRuR+xg2EYxZqrecHBSnpdEoQ7G+uGxQKGgs/t6o1zIwu383rf
KHwGGpkLvVlPxfsfbNd5hfiA8Ek/+IsymqD5pTyp+hVl7QH+aBIkWEp5A89l3J0S
KDnWncSC/sMKzNtaCxbc59k2ngWFfhnnx4/G5CVTchzyEbemPhdX1jd5+4/rOewx
4LMVPDRCOvwGh5d6ZugZ6TvAB6lQlL++ZuoDLn6sLX09C/WyU59wa9xAGaGC6TyI
fnZ+FphFSVXG8FFO5powql7mu0HtgIdnFiz6R6aL/FECsqxTj/CWL2mAHYSfG/sZ
ZZt9a82PXnzIHnzHFjFx5dbqyMV37DZQYNiuw8nO3z4cBXKLrE5jaygesy4kNrUV
YO9wbuo78wYp8agw5nist0BTS+/jk7mlfihnp0sckaxr1+Afz1BArrJWjSSgs1VC
08XA3xcfGnlNKjhSZbTSQ1W1AqFFGQCEMvFlzMAeZr+K58QjTmKLigcxN5OgmfVT
hyuXI1/nOYupfZ0V3sTakjDCIosgQAK6iW2Uyt/J7IgKsssAANxNgnftTs3XzfsZ
Q/EQJAFqTBVrxv+bo4+yylsY+lHE+wIl30RrlMW72R8Ptt6nyyCZjjTaIfvhRAbB
1U/1RS8GhfjZPg1mc6Xh95n05DRDITViL+L2176mxULb7OpuItZ/8kt4BdHmafU5
+Xs3rHh5H3IFl78ahLql9JReyzPyTvopbd6xCVsivA18VPajm7Z9JKHzkIgg4H9B
JGQ1/BW5XK1MNg3yJ1FEICdnqokVOTnnJrWbtrqlcAGENda2dyzRZZUSwaB611Yo
Cva3XAp0fguvXxsjqlSZwUbyJ5Gy+ky0/uOTPkIwVCIErXft2JJkuBempnP17jEJ
6pyFPgUugnvPA6wDVDqeKbJZbtQC9HuF8HrzrQnvogB4j60Yf9+K4dxpDOKaa/hf
UlFZpOJB+Z1IQKtP+PGiodRaHyARQYQBfw9FRj4mGtxugZJ5ICOAqoBMy0Za0FmK
vuZfce9TaQtPLQheAxC5ljJXRa7ELY13Gn8XYY+Lk9BKZVjV1EPx+lgIHrt1H0uX
JGJw55fHvpAyA8M/t4UdYaio9oPxJXffsZ5J6iL0m0hv2swp8o6spISTeK5jkpj5
x4lBPwIWqh1XY7oepuSQNsUbfs/421By2ms+DT1XdjdFgD3IbtoQph8CMTeWyPWe
4LEJQemm8M2mAaHedTdgmZjMMesbyBvTReOqMWVZvOJLSf33lPSB3q0iD4SQYrkt
AqxEVeE7YswcHH+hZ7q5VK1Vre6YMosouwjlJkfgmwAIM/J26JPSO9f7LvyAacic
BfR9AIdhjY7aD8Da48jdUjAfDXS50FQfUvuV4riinkAiNIWETTruvdQBPQTL7UF/
bRjoO19vZi78E3dE47dIi35Gp6Q6q8C0wi3UDrpUBSS3zJKWmG9qQ2vu5X/by5tJ
pU8nBciXfNBchn8urb72ErZ65cOMDs3ND/6zjCNTziezzKbd9595r31IhZhEqgGz
CT5asDnvSNN4G8rXX6f5h1g+A4ru8GGX3E4YyQueFvOMyZrmwWuvw5d5ASyehz7j
yz6oKPkXxaLavtZmuscJm3Ak7BOewdJcbCT3uZ356S/ZGdHykZ9cdBD07QMwojXe
T+i9ONtblg1SlT+GIBEJWKQ7F38256KaOqZtrJXrkxR6XnrvNPg58pC+MyZplKbI
n11JKnuW87FSnpiowgLKVNeRWvdxbBnCtzGHaHLHP5VCRVG7StC6nTG17ofv+t21
OHZq11lGFlDnbidlQCAz8ag8pZSjv88PQaUIMtL8c9Sk5yXp0kDScsdYA2B72x1r
yIeYOOlqzwjDM+J/w+IUZzF2M3w/S1NTVzFLnEdamZ2t0/8mLO1v5rXUlJy/tzqW
d6zv3TitPZ1tcJGbUWGHmYK4Tt7E6ncVHEoJ3eFn+uJY1ufA+yrdvFoMzHKNwA1b
m3bNXNiKljWw5EIT4vmJfO9PtrtlF0JOgG1rt2xjYRmQJ5BurZtU/sM86VYWKYOT
vLDRIP2QCFmLKVXzKATj6hutSg6Ea3dYo6fUAZnb2awEGXpFocBWk4RgmS2W2bA6
K5QReCuIt41WhoGEmqBBP87u0DO3eDjNxgPxDluezudNGIf/l36ln1gPVCW/b5z0
SF15T/7i3ejxs6ZlcnW2POhbTORaupg9Fwc7kfRzaI/mlXCgLNRJXDfYKmo1LfNe
1TEgtdbgmifK2koCYeV7eCJjhRO6wMuDee7ZoDe7KORAWnb4KJqkg1zSTjU7Hx1d
A1S69B9EYN9PyqsyNlMnFaqe3Zpt9thbexX2PhPO50S3ifj3zFcfy5aYdHAT95ZF
jrDSUnjeQr8BFodk1NwCzo/mFUc7lECvfCo0tfP4dvUB0/io/JMzqxPrKPlzNhyu
IloukPDi44Uv8rbwlD+2pXKh1bP4nW3J5z0bsykbHOpUV09x2dJLBLOnnpeHGnyR
epIe//XuVWFZ5+Qpf2W1XuO5fh/iE+nEUrzgY7azReTkhPbZxZ+T9kzVni56hJ6q
v14O3Q3LWdpaq+IqB97+2/flaL+uzt6w9BabdAHk5tNf6oC5MtXShNr34gJ3DNCm
7rGHkK+t6xc6YRIxBHntT0RrK2UVFbpf5Cm0wSNFJJniczudpZmCBNxF1dTLAZPq
uERqznaQWqzfig8KgRzvVaTIRTWXTF4tohyAm896GVstAoLDI0z/Oaji+OS2jJEV
0PN+Yy/+5RROzHtRdKCDynsbuodv9+wj72lxZtCOQQii3QuVPkYoxnWQxb2KoAb0
gj2fZgOHfHZaa8lfyvEhWPOxIqvVmCnz7qoqPlTeEnp3TC0KZuTF11Mq90wDQSnF
Gkr2iVixopB0tTzXx2Qnx8xSsUlIERdjY4NHu8Ak78NgW58N1UbviII9w4nWLfHA
C+gYxOQWBDezA2UWnhHxt13E/ATigyD983zxbbBFI/Y1Lche1qq0JqaLtbbq4eoH
RshO6eRg5/m+WXX08R6INb556pg08uX9QaVXTwtppZ/oaK3ZHOj7oNzvydC9gXmc
LwptvyeHRCamQLUvNX3NRXGC+fH9ZTjKsqoUis7B5ibGyA0MdFsgN8yuC1ZeQRLM
FrXIHtX8koBwtSXyGFvDNYiMDuBalrQRf/smnHu7Ilb1kLNvA0XWjrB50A9CzfWl
hn2ULh6fgLidYe01DnZx4fhT1FZSTWEcIp5K9yU2ER3Qn24LSqB0r4nBLGzwKUnD
UP3ZdKF9NHSr5nikhPCzNHnxc92FnQO7vigVO1nB1s8NU0RkSpFPFewBX33NDTiW
6OC6b9aanIeijqIBRk0IYCHAxz/yWBQ+tsf5c1dknpL07MboxJlGeTCeA09kx3Na
iziXQJIAsobuKpl+Nw6a2TF3/lm3vzZnH9KHzS/oxEdvKgCi0jmq8yxS+lp5HO/X
fAPBZqYdBDoMlIlfdEuyhH+GrPR8ZCKoNdiH4EAqKqAaX1m/yHqXKYdHE7910TP8
8fDrrDd1TFknV/jbTDUucMkpSfytt1SObpcchecBBWjHWEFHKyyCBAA1lQE4o3JC
hdwh69zCNEaI0r3PawffL9cv3EKjBvaMDLacl+iRk5bYYG19rg0yw7AzL9TA7zum
fx1f24deKOPh6dVY3W5y5/z9Wtuqn7Lmi3I6SO0/QETnB+hJaJkCwH8m+CPbRTlC
NNDAULGpQtNROIV8TD8mh+AqdIJN3B0MbbM5sIQciK+0t9xg9xEwSP4mjl4fMtj2
glbYdesjIqrLukk67qtNwcG7Ixe/d+om03n2pqu5CmhE6w/dTTcsq62+1zywb33V
AS9jx5UO1qVVRoLH4eW4HqkW/aCS+sGq5H5cDG9cVjqG93KU+dSKsCbr/x8nKNw1
OxW6gIa5EWerd9A1n5b3fHAcpZATA/XFKEOm9Uh/s6Y9dtlE6blff2uI5bb34ccw
dZUpunMEWMQ6kSzT9x8Lv2XtcmZlDXuJTqBtPY0ClJnoJHrwBWGmSxo2xnQCszaI
wZijf3hbiXUEFgXgOmRT8+nwduWEi9CmBIglwBEqi2+C7a2ZHGYjrRPardOdGOGf
M9N773CvE+UOR7eqw6zE/fAlzCjX6hQ8VZiaOhK6BjBY1bpt9d0N+pv8Q98sTheO
K5G/1vdzwuSASE2ZgMlWP9i0qg+Fiti3+/JR0GLy93ZTlutk7ExRlfCZb5vxIaxv
O/NSZpBFV3KQ/i1wkQ91cdt+/h/ZOAtleGUSfOZbvI0XeFaThJXtOQuFA2rQ9sdr
n59FVO3UFwstzxE+DlJ7zmC932IAeCumgTOgnMTZuwE45bCbv0uB8RIvQ0uzdb7K
a1QfR+3oibGIc+OcJoDqB5R8/4SA6kag0E/QbNpbZn/AZHizXSWc3S3hlz4ZCajw
Pi1h3BhtJIc7NFbJ3QMWatRf+sNncQtr4iSoagyt2uztldLND9rv1zGYvjFlp/8q
28EV98A2w+dm+I1u1k+LWwT3Zjkl0xUxC6ftUScSXAXBEuAswNEhV8ji/xe3qqu2
Tn+cioUrH/K4N1kBbHqdxtSx6sFpvEkDVb2QPlX3PtVkjDjLKpQ/KibmaOwMoBGj
tIeuOPkcLwAPpsBCIdg+j5UsZcVT9WbZUSXMzWB66lbF3ezd+7KxpQAz1obrTQU3
xAdNk+4h3CLowsftgeNHKe+HycyTxWvc66pmFREoST9y/ez/OfJAXotEvhHGhaKz
QPKcmJYLRKhmBbVEVbLylq9AmGvuMN7mXUizXa/kDshrn2mMudvf3VMw6GA8e6kP
WBHBCvkx69Axt8zQFtlrBE1VNKrg07+Yugo/huJSTHv6Ti/LbIB0VaRkkxmmJRSJ
vbzIpBg7t1JNNDDB4NrKWqA9z+SdSMctloCAgvA7YeyAZrjWjuYlYfj0Q16cKeCR
OjIrOfoTh6X77fkX0qnsfh+LeSY809GDKNAdslBbxxAg4az76eWvZbScq4SuYm8F
JkzXWP4E7oYl+5UaOxQMnKXOzXB/DC7nB9sBpbBpoyaXtidV8frjGekmrcuJf2Bi
scFQ/P6CkSJF+XPlzu9jWburZiM9IOYK8xrAFNwAIfvBWuVzJt5m093AGyacigsU
r8VfRtSMSTZ/JTaqaM/E1ykeWfgDLX7nXmnKGA9j+WxE6HiyrAMwBoz8D+LCAZq8
uBtHZYt9IUMApv4tSUM2ZAYYOaw7Rom/sHQhUpLhSAvlBRGzFh0P90eRISe3ckp+
7/xIAjLTEC9d8/F40cwdYOvrekD0A4495DFOtelYLyvjVGF5ZxiCuCLbc6IxR+/w
a9Rq79L1MRQEeDASyJlVRGKvFS4MDAQrLd+SENT4wW1yXoCzEcBmSWUKuWy+VpDt
HgpdNoEQnhHJd7OXfhiqqkamOhiZuLfJj3XWU9MSov6VF1r9RJ7YMuN6Lr3c3Eky
h8ioeNfZVYaC0VQdLN/5UHMbxQeIFX5441L1ILD+RegX3ltGWe+8rXx30cHeQ7L1
o8BpBKecTqlpv73W5BbCTX9jS68vKT0/Zq0iokbNp+VDjJZUq0sUrzzLPqw+wIpK
6t3VOsx36iQ1FlI46lQcAd1nYYYgyR55wA9NFXwUmN7GTkPZTiLsCrnvNYceInCm
p57UfDexaYwwQABVyFyKEl09MmKQIYxJh9Z9442dH+LW/d1pHQCnSOXWesTtkKmn
j+y14odhueOydHs5NnvRYbJJxKHZ78qd6IeEQXSCmvPaDDQ0lOPgMOVxTDEbJBaY
XfyV1K0kOnwE2prUkpmRsu3QzHQVQjIuIVpgVuP4hpMxnynbibYew/jzf1KlnzT9
xMwZlKFr37JEdNsiYy0Yhnb41A7EzhLe8+HNy47GU/Dlek0NTSTCASuJJzpDYrVM
AR5oWS7Cj4f/PahM+TOrDbQ98o0z2M9LhEysFNAf6VH+9qKRo+9JIthuVkG3zTU3
d4eMAl9xxn4ElST5l7Eq6d7KtI210ZM4AtLnNf4HnOvnaBERE2RFxMQCkrHybGI9
Y8T/5wLqGF0RmV14U+RcwrYq8L7RQuKHGIejpcQLQ2tDS0F0Add3ZrGyRI+D1Wrf
jKmhUbU1VkCIHrN7MsrnkNhwmhDGjO2E3fkI043k1y0K4KV1gdwiL27lt43/SZh7
XMyzfCTr96F17FJ9rfUPljOeBW4Q1nQ5ZOWVinWrtRTjSWbewKTfAfZJLMlb8DWa
VPQosGYF0rBKV50M44Jquk7h6kbmRIKqm7RGVDal9B2Ibe66vmNNYS18MnXyus8B
Ia8GsCi7eDuxiNerDFQ86eK8j6P5zVowHtcgX36kPP0arTBYLCkSoam7bEMr8CCp
cpg4tTgc9TnTPYlKftOCYfj61MixN32afTK3pTd2dAASAphEqJ1hy68EAG9MVtSd
qMGyjOs1gVlQzfo50a7vBRP4+IKepzeiCMPIrs7trrPU7HYkvCkyd2BhkdYBF0aS
beu3uN6D05vKkSWdWeBXU7VwDA5xHGdTk8LPaRe8mv8v+I471dTAbOl20/J176Mo
6jQmMnwOyR/VV1ELL4ywSP8SXvdFV4pxoAIwZ28yLBCUuMrD/itj1mc5h6ol58Rv
OUE+fn8Vh4xT5yeqb36ODs1ue7TbVHdOxNb49IrVCrUl4yag0Q5CIKK91wYqXZ5y
SFsZ9OiC3FrMzSSkVyH3tVmvJwn9GRRUFLHMOfb7VezqKgQhpLNcD+BGvagdB2lW
CQdSeBvtA1jO/td1mGv3+8x6apzQerLKjLWXchSWTP/ZGUNkRbfLaAzND/QN/AnN
o0X89ewWCTtHYMNDi6zl6FGHgdoFmrbKHX0/HeP+NRSRVlHytRbP1c90Fo9iybXY
+DrotsonTdoXgxqmkEw6XdzHm39hC3R342wxLqnTpPik6QACIsTfAkQy5G/lS/tt
RAcHucmPVdn/Ub9P24xIPDAWUCzwVyiXV66Spbmr25917i5P996tg/xnjEAb6T7I
DDjyOUgevMM4/qCnmkBwcGgMFUf5x4N3glwhFMlB6L/bbl6L4KnxzetgZXxyBeVr
6qpSVj+hfbmQ+y5sxfOtw75UiHJrA/KjumzbRSk6w138WisXImezuzob67CqXqz1
3lmNeYom9Gg8OeGFseMuPHqVwq0k+e0xWZK5ehcnoc5CLe/wnXBUE0qhBduv/OJ6
+0xWXkBKbPARw4j8gI3QVVMO/pU0wZTIuP7zBm7R2xAM6UFW+CJyx1IuAz0duT6X
b6dCWrlj+IGvwBfhUYepYbT7gKOuVnHDsI5UyBevr638tAIwBeoCi8eyliDIlfBF
YSyVOcAwAwsGEIaQs+os+1lxCgV82d9zy7lupt3cE5fvJcDpscFtS1pCmiZod+3P
d6VbATYlZtN08H4BFyQHp9svfg9w+YcBkgM7+0EV5AvsegixcAgrEOg7Phm6RbAS
3NLa2J9jQ1CzLR+B+w123jMOb8mniD/OhywAbO9+25XtPHEsDkjwFkIjRXf+px4v
INz3SUGj7uvV4oxYzXMKBXhzUJmXJK31JgYbdv+HOtwPsng87P8CDuiPHSQzhxGz
QBz2uowTglHKrlsllPvVRVnpgTeZVf3iIpNa+UiFwwm6rSDy69HxkGTd6taJahIF
TLlXYGb+5A/TaYuorNMbgc7n01hAjteHwU1JBJRJxgOsGYWh9VidNhVG/JplbYzd
4ThDnpX9/JFFSiR8Rl6xp5IeyVb6zYM7Etm3Py6L3sr95yvrFEzbDgpZiQP2WV1i
WQ2iTbURdGzRmqddwCtU5nrlTH6PRyfXczutUgU2tLasL3wbA86/pgObHXUav4j7
ym4MbTUvKHAtbQlt6m/ChwbNQjjPAmrXDfL8pUE39GzaEWE2GjliWei3nJVWgaom
8u7Z54PXGXghA/TB5BsvKlQS/n8SLkWGh9LJIptosIGvp4lvcy41SulQ6rLBXwRX
p0WU78uuv3lfwdlFy5Ezp1+pssUhwKyuDyPXEkqaj5RfDB3QQK2kmj6iYWk4mKOV
3wmDd0hIN7cajZ9jiZ7LE8sJGJHRVjHYSpYU9UNhKUMNz1jMBjsNENmFsZJeHJWO
MAmP+jixu9egtp9zghP3oSQmpZgiqKY9femDjI4YzdcA9/t3BfOkurs5Ybudc2lG
M7LtfvNVXwZE4KuHRUf9fraqF6SK8Cm/bA+QtR1Qyli6AtWTko/bdgWCkXxxDqUf
Zo9nk6MWGWRNJI9vqpbBuwr1gdrKt0tEiggfrscER/YrSpaMdv+xPiNrmtM2pLp1
7uAaLe2HEgL9LfSj0eT6DFzS+vfcyj1OzK78TPy8M1xSCQetEvNujTYlY27JF5+c
miIIouOohaoEBQKFhXmhuCbdDyzcv3FbETgtNXyHJ5AubFpjzRbLL0LvcH5L6Na6
tIOW1Ow/M6z+VzK5vIX7gKOQjhTcgxAAR1p7FcmFW3FdhL4d0HvPU9pwWEnil3/h
iLlVsnUdf6S4q2tX6dedHExD2NPW1RJy7muqGLmxhEokpbXtaZMircqhY6kcTzcX
PwjXtwD8sRRQ3OKYozO91sZO1MQtcSFb/d9oT1rjm8Gvm0c0620mSKC8TPr358FE
/C5Fg9p1qtaTSRDZcLmNxSO3Qc4iQ/LutGIXkkeprNTP9nsthAo4hg6241IQZuAG
Xz+L2FaQUIhz4ICm9QGmSNFNbfXTZ7k/xGlFEhu9LiMlQ1WTjv741zktEt5oz9FR
UeHjvxOYGRAUC9VBy5uZTy+/yVJvHutknyDKHUVH4hefDs/oLsCwjrgyfH8RTxAD
SsANniauD29EYftjWqhYPctj8QpCw4GPaG5epX7WCO5G4Ohm5bpZ+/OOVMC5Emzh
RSnAkPFXRJRKD/lbDh6TOGJcWZiRzsvMn2H0AZC+8jLmAMfkK8ziZD0tmPvFs8ex
fMucBYmI94RJ9y++wn6r64B41JxYPeXP0KZRn8LbK0mjnZaAAZOxsKpHaZVSmqSX
BY1U6zTXw0v0++PjScQd4NQQxkUTPsSt6bHPeljW0sv5CtpxwJ1+AzK6qXUBVWri
CBgLL5NO6qydZLtKUksVci1hXhipbm4EwvOJ7gDDUIkfXjU6ltVxXOF30OhVpOXe
3OLPRLjfU2evf97uJ+fTG+rdaBPqDrWJU9zPmf9mmnzVWwKMqEorWPElhX2TjqBo
WWD7SUbZcxqwufTdT++DmWlmZnji94ir7pJfzPRKcOoU3Z4zjZH39ANtCRwFi6YP
qKv8bJPA8b4FknHeier8ra8uA379QMTJ60S3JYPtH1R4gWtvCicgscfeBcGKjhzC
LKnsKv4WBE2pBq0cA5XHdIWrt6UdNGbiFXKHmfiNuUrtgI2ts50FcOqEcUzM93iw
hikiLdkcH1ngFL2HZkEeRoTDM7yLap6vAd2/5RO2Kr4L6SDaNX9GXGRTlV1D6Glo
VQoZR/yflugIO2vft8CWnODMLgxIsdEFeKJRHm6bTi3hESniYRiDXW/Jp89YSMKW
bcAk/imJ4jhu5U8acm0H3qjJ3JOFKg3RaPCDs8SLIuXAcueSZXE+2uDmG1IUGITg
Do3rF4zlVVSk+fOo25SVbKkpbUS2pBdwRCF13V6VqyEw92XrVp1xxPrbCIsDx337
X4ha/nUiZmHuqWq3w0V7OjsAFfhA67t4qjkl02d+VnoHeA7fn8LRL6kAsIrG6+fy
N2SzXy8wCG5TRPVPF717Z7VjNiR2noJMLK8lgzS6ZFN3w9MNfDS7B+Ph7W/Dmanf
hPu9oA9lWEezlXfczTI7vsPYhnvDY7dJKq5PgLhc2hX00vyIIIv+XFirs8bU8u3f
4jvo8wyK1Bq0iDNMim2oKftD6pGRPfPAL2IPbf9ejbdO36+6iy5JntjFIrOIrOXD
LN+eSPKiME9dErSdmnpJkL9GLQAJ1AfXlMFJcI55fK7DlIyg5SPVg5NlGkTeo003
rFEZLoUppvl9uS0mEMuTuRuE9HJwP/vAhxBtkiVN9co6JQ0LJj5TRWJ0/JpOJ2WR
d3DGi2nyRpGPBU8Jn0qmJHLbYvxyXnmAVRhT3NnzJCDa/D6xFPHPFADNUJwiZ78X
U1WJY5237Nitw4LfUxjnhGthzm3XdcBINQOqEz39gPaEoAistCfg9l3oRtnuqCHI
8qlC0RXU6/0xyP2oY1fHZcvJooVA0vIRJmztnbSNK4wojSuQJ8L0zwadIgYcWDbD
DSZeR7c4gtlkJzCk+9vIGDq+ricAcBeQa7eVlCIOvpPoo8F6DKnWUH7alWZxoH5V
2PzbKfXJpeVVn0c1tOR2EaJ9m0M/JuNwMq3IoKpRwmL9DxFKmyppNnXfmI9TzyRE
/BaT/lpEi+oIUDOuicD2D0YcouXKTa+QKRLv+L3h28krL636r0yLlQMWZyERnBPL
nEk410PLk1w0imMTfSsIKiEGJsvdAkVxq7f1zF6svxM34Jh/UPdZzGGcRw9LLk6j
YuloJIIXBU+f8jciIQ1K4Cy/j3dRWWtUQsdiHI5nc753x3S/KOa/xLX2G2AckC4T
35GU+4OfoygZBI2dee8E4YAP8J81s12c+QiZphpDJjNChoz6BPPHMGU2wDwAAOIn
DRlbIhj8MUxZGbn2YEY2tHGX+etTvurldyvDCZ1O6uC6KMPeTs2YogQ1NzLKY+0A
ekGNJU26d3UBnvgDZ4xK/GoPOyLckGFr5CS6v8k3AyGwNEzwrukSsTCOmppUj9Av
Ki5BAPoZR8BPYPPz5t22cUpAtn/BMSSX/q1n7E4K/5uwFwnTjvo7p9ByZl//4EQE
rFUp/jP3tRL4rq45ZmjEGs4yvw69u8wqJf0X+h4CXsjT8NFTiDg08cX8Kd/IdWAg
lCUpADiNBUhWRE4xDV/gpSaVwkTrGoKiJkSOUMu/EarBqq3eWwzP3pf/aq3Lalce
nw3W2Zw7DrgX6Oza9UfgOytm54IOYvgX8ucg3kMmT1UD0+vqBcU2WxO5RbXfbbQY
eYJ1raDAMZapxIdZb/8cMNRlIGsWWkAdlkrAZLnYeNxd6TzPSs0r3k2nE4Yn7+KO
duS9YecCmTkil5rmGw0SXdSZhEddJuBzhXMDameyoztJm0uJpmXeRBd4zWQ7sucE
UwJYWPnXYB4cBx3nUjEYRtFUzmZLteBb4klRnDpDb9ppMfImdghS3LpU7ffYc2uO
+IW8r6IqIsQcU7p4y4qr2MVYUp9VKgY4u2zGdtTkhRwtg+xu5SkCfdJdKFegT2te
MucXKzFFCCyspkAoT9sfSuN0Yeqs65x5uEGQ0U/qrNFwbqAWKwU/Va12Fxkz5+Yn
VNtk7hio+VuBZD/rp4iyaSMVcTR/ixhZhBsqX8+Roj4RwQn/S1MKuU7aMm/nOp5m
Xd6MFc5kRDe6gkyUcpmq8SbJKg8+7cxk672nl3U2lL0IU3xuTEhWxrQxDr3pTsIO
AJafzVPuIUT8bs23tGabAW0zyEomeQQgQmYF4J8NGzBFkfPIvVOX9z4MpzTUVF1g
CqJbpF0lWRAHdhyJ6mORludJ9eHHt9ZRIQRwuVsOoVrBDWjgdkynhT/f8yFcj6pi
M1NLQNIkOELQQUv0AIh+fpa7ukTmiZIixKyWVjQvNj8Khx6zH+7Nht90VC9cQa6A
KYHAIsSVj+lTlHfXGC8kD7vDVCG13FTP7TPBiZrt8OyAL/TqtV5YUsK3ayZzlG2M
eupCSfWZyDQpGllmA6Lzd8NRivgT89jvtgga227cOeSpFaoHTICvqly6YvHEvupB
3HJspzIIqNUqfd8QQ5rVeYE87D6MAmTnGC+EbwKe3BSmJdyy3MwPNXozVz4IxmTA
56u+RbrKIxwoE0/Xt+tQ7E3QzDbeh5FAovZ7jYfZzZEDBscCwbuOKeKedTeT8xiO
Vph38Yl2AXD0ZhMgQAejQSOpSBaw2t5i0zseDIxrn0DenX/oYWRanxJfR+XRiIin
mWQ+YULFxe88Uwn+Xt7Dx4PL9uL/bGoQvVwfnXlp7W5JqqLRrhb39o7GcpUvOCZi
iU33Tpu0Y0Z1F5LbdAi8pSM19fmNY2Zf8RaLHizQYznziTnh2GA9qgCR0YXsZq5J
llb8ApiorMTBhn9/EjPI37bbTmmoBhnyBWI7qkCbQHYAe3+SeLMmiU3yK1SaECFL
dbVQa+4s9j67QGsSjxYFKhJyJfumKvJUN9ShybB5dcFHEcBCoR0fNO+f+Jndcucb
a8Hxf7N6EqLpIABK89Cx9+Syb+MZGa43+WAww2NdwVDb3/r66wRrUNoAJf9Qev+N
bBbS331O4i4fPuw23KtPyI4X3IPWm1nnhdTkLMN1M0Hc+p/phsOQvN7WayLVplEO
7rrQgGxWYNrrKj3siSqeYmMVuEXtJ4xkSwjqb5McXtnLQDQ61vpIMnoxnD/gIc1R
mw33wrFe73Pp56i2iC4Q2ch1JjjB3yD7pVfr/hlTDzOd37vFjZihVL5q3SpKZmeb
EoAoogF1Z8BHr8jpFvYFyY2EFnC4UQpBOBORzpL/Vz3GZ8KmLBoV+w13UM9ILJsZ
h2fYm1k6aRryITuh430m+817lsTX0HPqu+t2gDQFrIsYDF0oWcGKIAyDN2Zppb4Y
eYaBv9xLE7YGfg4N5aNbeA2MGWEEQt8Pjst0W/JRwqBROd9jAG3kocLn6l/+GeP8
VFBZNfjabnxuJ00g/7aPwBpzq9S29Jyg8tulOwTTwTzai+olLkAyc/OTfiwQKJqH
naEN9k+kqPH7p30JjIwFOi6lwhErcn6NmmK1zSaLuE5XunB6R58KVQoSACkj+/yk
3ZORX/EX+ybqP6zr9d/AJgZXJRtKwjOw/FByFvT4InyXjLBxBIWT7/hl7QKIFHNg
UaB0hMo94NBJrdZKlayf6QesHeJ1U8eZDDsSfMwamQq3O6FT0Mfa/rYW7r1rrS5+
jE1ouZ8G4GCqcWBS4UgVZXKjl3sW1ip5sB7n3gtxZHJcTP+JT4zd6KvPbFnJiIpm
uxxAYVZ//uSviOEZIwmj2m4E3z+4TbLIyhoMzxqIYr6+jOOIs0yp20blFBeoN1Xa
RpUHlfTuaXDDQjEwEK7Egtkl5nr+j3a/kTYvU2TKBPeRjdqtiolXAuLdfJX5O0gk
D7zUONjSUQrIS98UaMKHkxlz77wnkS9Rv44D4+OP9sp+JdPO1kHC76wNcraOH5w8
Qx+VsLFX+qMmoRTN1zIf/hXj/U/ZW/svaW00qXrXzY77Mhe2eAMY0ZjF3w+jbD8w
wGK9MWNDtOm1mtIGfo91RE6ovs2FIZuVArEsfmRLhNEBIAlqBPRtjkL8JVLJxEJP
NQ/K0/UWm3asODZTkX6MASK9J0IKoMPynUFHI3h+mbRQn8prCFL1/l224+bO31YU
+EAiRzDJqmPWIXpnjbSGWXYHjZPbd3VCznxbvpdpk66IB6EFXka2aurMDeyRaxHx
1K/GGEiyq/Zy+upZAHMPLRWcv4+LNNn1xyJ5YNdJWBXk8dcpD2gIrmqblx6weBVn
ifpjo0902b+shF2YXr8dP002MgwrJ7uMHU6hpKPTnOY04qY2mNrDl4C8J78uK/4U
kphLRPTh2AVZ6lwz0t9hS5e41WOa5z/0xo+ubAafJZBu3m0vVcTN/BFG1ubOYaLq
WEPpue8MaixaMvpcGtGPNuQXyvD+CP9Q8V7/o2i9WCBITM4Gqo0zZYkR5qsTyEnB
U4WrjT/3LqT3ELDvJCOLUMIUGgXL/+H1EgSLmOSKApHldDg/yJ8wDSyeSZUF55a3
CSr/u2f48DsEz5hT7nnkAmtduKTLyqVf97M4RJvwfU5lFPH9Q/kGJvXzjBe6g/JI
RZcSe7oG3B/jisuzUqLXjDTHovUIFXTBBrQ7OPyVoNGbFvNYEz7uGCudonSZATN1
K5fwU5+FuZXTfNObJcgc4S4Q1AIUvGGdesMIGX3onXuaFiIsKqy007f9gB2RMZir
YqI4qqJngAfKkt/eYgtn380dvpbg5j8NENfDRLo3K+/oxqmYynHrcBVZPp0H9U3Y
Bi+FrE9ZwJt9QwKQlu5xOki66AhxUt3srmnfphxkFIdWjD6ZjEfGeuAbiuPSADPv
C8qOpDguHeWDwGurBBXMs9uK6IG89JLZP91VwV/1bSL5+Ma3FqXZDg6ymfDT1c34
yPaMfK0Qa+LgFv+SEI+fEGZB8LxbDDSPIIEO3xNJo/k2YNVUr87VzA1LGJn7T3Lp
YhyXXy49SJN9elbJ2ERBGpzex4WKL1vxPFWESHHEcHPU1n6y6kTQ/SMiESFQ5Mk0
YC2HfZ5wjTqty3ZtAW0P7t8Ylli4qys5iSxDXgGyPi3mZLPZEwwIKbtjBZNg8Kg2
tfudVqW+LKPhO6Ed9Z2kxyGz287cGtOhbIGd8oySjzGiaEkoZsTXdJCFJizOzSRJ
3bl56spG3Nq5VA15M95qKO6NXN27Ly1s/6KTS9Kc/ovj9xGhf7hib4umCYQppUb3
SRO9RLlW0xzHAWVWJ172mmjNnBMRejpUYxPwHscYZQV8sxC084gTa9kf7k/5Gk7E
609iG+YvG2Ux61sA6mqh2e5cyv3JoAH+eEDvtyfx32GlR/ZD7WSvWFovVLS5VLwA
+4/aOkAdUoxzAFB5G0HKtAoSbfrHzTXBbLh7I1szQt4E8k/9KZm7nl/QlAwrKVuv
dit94LdBiWXj3IEWA9FHocS1s29CWo5qqqMIeAmj/nOLKSiuke8BijpVKwnhYIX+
75AR4YYuH7QL/ShaCGrJKsotVDZ2cdoCbH5HFiu9wnahxG1h/3jkn5mwEk1lg14c
J3Q7Tt9IONcz4Qp02WqfXX2Dty5Uw8knJfrYVzwvLA5qJxdG1pkdhNxIbBwYU845
jMqdeyMHUqRmqsvKET3PVDgbIrHEavke9n+12WgdXjigqiooa/D32Bq1Izp+wOGV
kvFViYmBxaxGVClWbyEB9Jz5/plhCz11QMJA5bMZGqJnqnwquwc2ihLzMHNqxz/g
JE2AbwEkcIq5ayhTX9HsdszufUaO3Ap+1mHZ1ZlGVxkeZ2MN0QQwoXkZE6npEsFz
k0uPqZV7U2njVveaBMfSjKnZJx0cmWCBWe47FDiJMibvvDYjfbrQIWYJD3o02hj6
WbCR9vv8R/ul9upQA9w5IUgxJ2zczXdj+90VuGKP5Rh8Dxe/cYLrmMWtMvnO9HqZ
UxG2eajMNPfKlsUQl7oZEYd6PHf6AJmbiiixJ8OLiv+YOkRESKY4lrwCJdS2Ib7n
3y2mnMuwC4D5yvXRJ2pGOvyPKjgGfayt2TSOTSGxDco8jftHnGU1GaZjgmVg+SJQ
AKhT54N1JjB+uVGca5PzO5jtWbQWVRX/GoBBvJDAZxLKwY18MqRUkCmjjAmv74PN
AZloR4S3I3mIjrWFby+BEh/nZTJcUUHo9IeMI8Bg7MCEm8XOKVpEG8VEQtbb3b7a
ncg0E8LMH1whTgpMN7PBcXmUEt6vlbekSTR4sxhYloMDrkniDcrDWt9+wvzxV9/M
hXJTBJBYJ75spXS+KHs2gS3LRLUuxdhHMD8z1SnWCSCLd+pgNxQvNK3oZPI9Ph49
4YmSZ28ZOwOEs2tS6BKGV4Nv8mmI8mRh2P8cp0u3G71ZAbqUtRjHeLu6NzsJwj4t
RdB908Rnu0opt4ehULEfLWz3ShQZeNgMKgqvLPCgFIjAsMzVRBT4Pordxsc0Txaf
0W7nLK17BZenaR3l0PWThDAOJV23I0/qpH3O6Zv/HsQ0nw4oIEMpdDx0c2EfkCSr
KclaukbnETZOSxMW2xBL7AS7smh4u3aEDffNoUVbNnhY153w5TFR89RHsV2sTTFi
DbhdhnE3V7iraXPn4zGyxZzUUitOPfc7exTvzI3FioJKm9bLEjIwu/9xAezcTq9H
6ZWhMU/smgi6hAF2vUcj0yasYXPfd/hCvsgYku7Ac0jI/bdUIdmYQxleGKogyoOa
bvstzCLV3KFi3cO03xc4MMSBHBGxEvo3dXCCmrZQJoN6JeKJznJjmMizRXJCtucP
nqznLW9z9f4FY+nU7e9RwjRoxE7CRKHthb7i3K7BhOIV3l10OMfZV7afZsuNJUKC
FmAtzxWOa40X1Bs9XFRtALSYXLjlhha9elkRy+7QM3a9YQzxEWYXKEwyztnrxlvL
r/6GuiIB3p2npkFbhq8QnBW5oj8wEyC8EpuAJbM+ld08tabEfiGv/mKMwxtCstU9
RL0ehXHpCi514YzEAzRTUzFlpN5AqZkeJXuWKpq2BUzdFNGyxc6P20LAp8JJztM0
+NqncXvshmoeQ46MPDdR0Gt1jO/+YjFUvrwpnkbLsg+qze77kfkhmvEosNrO7l9d
93hcJlu1yNGPwFNkAGNaDEbai0h07YskFGCl/NlI5a5ZyQEV/kHMLStaCQ6aYn6n
1DlwIWkxBduTQpsf/xTz9gE2zEkFDJjLqDKgitViBvah9DlIWvvt4vhRLC52pudf
ZTQjDLBQ+/4ctB8DsI3iAk0Om817xZ9GcPzdTVvdaRGvY2ZQAOaRQuqqm7yJbxWI
OoUl7mPQglsGe3k68BKfeEtkT19166tr7nj+55VQ4Fhkjw+BfhbwYDHYHp7pULBG
u2W3FKAImPE0dn/5GwLZzFkzmA1PMgNphxP5mAn1VDOekjGJaKFQyDxdGmVWDvTp
QbD9CgjrIBe01HilybBHDnn+bSE9Kg3DqRlzMaXVHBRv57xFQL9/iEnxluDKWq09
eHdlUo4ydzJjtMAOD1Sx3P/sc1VWsWjIdzfbn391hqXvo3FHYSUIiyYJVRBt7hC1
snErliIjTSwFyZTiyb2ciQFnfkQkxxgE3P/uBg+V5upuDkx4Fc1iBC3Fiu79/tVg
ve4Zox2sz5acTKlHprLD0xhTV2oAd9ygNYWfXjd02kaE04z6YaKwObInnf7iVYua
MhcMr58+tx2e0YYaLEDKK4jL/7Q4oTUtIa1hCbsusNAWHxHxzdH2nHHwKUbgFHCj
vhhaVWxvL/8b/JdzdJeIMj+hvXr0BGYHCRCTISUnRYC7S7mO3SyU5U3SAV5Xj0aW
VBpM1e/J//MRNN0B5ivR3G3YVlg4g+PXHDz0Mh71uunfenBmpWNUfA6qO3bIlMQH
D5V9K8DsT2SGVEq+h3jXg8GGzD+X/nXg4LrJLa6aHBVEqxQ0Ycc0unR+srJVy+rr
iLB5aUtCTqXl8xhL96hRhVQCDk5EirafrG2HoIavaek5rGvJUpZ1/N1FwqGA9rjj
WjB/DaduT9Ypm4hOn/TA85GgRJanJ1/NdmlvO4KAJ7qUAcPu/VdTtZdcAWFKIxdp
v3YjTsR+SvQIk+4rmev9mr8368MkAvBKVP18/AJYsuesRnuezsVtdx9zjMPkmQ3H
w2TCTy30hImQWb7c5uxiO4qBcbSD3WgZihGoBC5+i0upNPl6J1jZlRTP1uesGmEv
XHLmuLdndlvFEdo4+y/Nd8MpIsXdhK+qcGGRY3VaulxV1i52OOy/ZCFWkulUW9gE
fR9f06r8X36UUEdRuZARLc+2+ZOLGjVq1K2L3yG/CjOXv3IoBujvP0/s1wYQr4Wu
W0O/aaaI4ngFkp/OXXoFegqx5Op1PGUgzVW+3/w9koHzlR//3a/OjRaUYvF9FJ4g
74kfVsMH5OWm3Mq6S+yNrI1mKebjjaHlCzFHoUuJW2c45+pkRG5b0S2zLggdPXzc
a76KwGZcvBVJl/+BGVBnQkehEJQELqrlkJopeF72X7eMsyQJ5swsfXefD1C1cUhf
XKJnki2rC/ZB/vosjPBCcaZDRx3e5GQtMiJ1KCwxlaVfc0jgBd4Qmqr8YQ1nV6iv
iAXM2zqAFSnOFnHbRWi98qj0pO9ruGZ5+IjpIAzRash1Chy3zJFm1IVILFu6G4p6
SG4QwrEBJFS1nvB9ScyxMBRfufQyVCLaRH0F0hXs6h4wbV40ID+8vJZbuYc1OwdZ
zSFIPSb0isXEQUqV6dl6zyeJg9sYai5bmX5BDkXra5eyO76DK4AJofYctwFk1re4
+uK1t6nbc0d/WkkOMeqfhdC7uIMNEtjn+ZcvhvFQ3Istn5ayoOk/bUW1iyu+CgQ9
hU8DbdOf81GBEfJWe5dsCCeTGazqpbnLZR4j46/mW5UDb0Admimv4cfpVKofgtDD
fEqRu5MwBt4Q58fIfaHUfFIyFdZ1pgJoRv773kM/+IK3J1g5RMQuzfnSHWqVA6KF
S30kBcMxakew1N2NNfKDFTXcA/b30u/6KRLTBiErglhM1di7YKVHFzdkf9Ufmeqt
IXkhAW+4SOJitNSh7gy8Wufhb/4Ga2y/izYM/LckPe3c6b/uKorlWJxy3yTMFnsT
8Vw15VsJ6g3moCmc2c6Tuh5SehBfGWW1uu+/q44Z/SucJuP3QNH0+wferd+XZUM3
Yv6dV8qQfNIrduW2xJJ1eZ97DT3GBZ6afHvE6qhEzgu5jY6rdJZmJSIMRdrAssi3
VQaofDRwQeffHtUxxnqx/Fvq/J3GzhfQ+cvWxnZa9GwEL/M9yyRvtpHmgTcReitb
O2RSw73gMYCCYa4xVwOJ0C09hIvBqHJpt6kGoO5d280+u/PjX2eaGpXbvLva6NPI
KiU7dUuViB5ktOvE9VoZI516orsj+e7QhAxASs3wLgN62vOxT2tmmZxptgWK8VJ/
Ty/fiLcpfUAcAJepXK7tclmjv9Az1mIKlPqWCAJrGxgYbzL9b8g+BGuy02pXY9ax
3lPa+Q3+qA3TQfDN+0lubzklEIelOiO9A20wzHu/JYeyS6W3jE3AindmSgwC1MNI
/g731I1lTmyDkgXP5jOs6pAikvqTsE8aMfiJRaIMhrb20J3UwWompYk4QJZC27gt
dn5N2+HHqFEa2TncxGulgySpGaII/OOG8ZExCesRWGMK19C6JuqffNtnOJouL562
BhhhOhCmD9q37xNWpjxn1VZZGBB+bwhgeOaAb/wiujhfuprdzx0fBhcSp8ek6bGD
bZWpA4Z50so1SVNfd6j+avGDXDtmHKt33gAIDWZQRmF6/8FsC5kJspZk9gvElidV
yt3VvgbT9NZvPY2nciyggl5wND0ohdRH4je8XACm4Mb7mx/wm3niDBc5bZqyiSzD
W+eRutHirgTEDuGxenPtZhdnpqM5xZcWBklVnLo2BB21eqBRxXsf8yKynHJsdNYr
IfPox/S8e6pf8Zy6Kg4rxUS0b2mnk0faZrqYZn9KiG1kQ9N4kFDwWLFdi25sjfCN
F/GrxajRxF3b+oQkGcJWaeHqBCS77ID2lXhaqjY7WMeuP+zdYgJAyvm5d4jhbCUe
RcU5FrLEjWhy7PpRyyIPrZ6PRNjL2pV3jwseiql0gUN15EONxoKSiFDJri4WJqoZ
2QvxjZJJBmYUcZNhRJoo3W5qW2tQsh0/r6jfjjPd5zH5HWoa27Q+57W8rDYZrYDx
9SS1PARDkwES1PXtzIX5zHEkyDy+Prhdarb0N0+E4MMb5TQ/Ui1vNTkBLwH1tPQW
1gb3t9xFO7tKbYWl1vAl/mwD82jaCGInJzynQTdiAtFjux2rzQtxWp4J1AHrDQx/
3Us4GbmqAg2lHwQwD6msDDndJbxpIsPPZTKg6N50xwOhi2kQ3eB3d8xpsOJqBKqM
QwVQoB4ht0X8Qn1n3cLYOgr1gY5NUFM5P3hkBLDIJDh87ZfrjMWFOQaPnq6aJb4t
d9TI896R/RYEJ7OCH+JUaKnOzePcAhjrEPbRB1F+d4C39VTwS6tu7fyna5ofuhvf
IXl/MxSWJyKaKVf11WgNR/aZ+bzRX0rh0n3jLj6sXiAli/8T6C/eVYjwdV+eyxW6
if4+BTMQrDyPIab/x3OiznLEBp1TBR82BzjvUWZfFLQzP4xrkYmHaQ9p0PKJfcvp
Zd7+peXG0JJoZesK7efFa0vW5ycgCs/rrMbzT6bPoZo4j3IZNSbyIyHEa+QFohWN
DbdAio0I2BftM/rwXHVJVqpz0DapobyulBVfN1HL5eE4ljKat7yxu+A/Slmchu1Q
rIBQnH74qAnA7p8meClMyYZJ/Kv1jBtZ34PYOuEKEp6KPIFfUVhfo05bHkghHQy8
35LEtEq4gPV7cNJuNJD86yrevmEXpSDVLJbG+swhvqSSEPQVmv0zFbqbu2UObMTV
1T2tUoTYo9HaQKgrG+iw4pwQR/TRyKAPD6AHoJKtUjw7oX5+tmh/00oCEmVPi3QM
Eh1Dg9q9AZr4cT8FIV5JAwIyMGTARyODS6r8yXaS/w8zitgIwIDFjpdSuqoPYqzH
U5n3IlpoAPd8KIVHZsDkk8XE7tyBbW1vF3ABRj8hHQPeqNRUwjIX/rxqxGJVyl7+
Wp2jf2PZk/G9NsX3e3FFMhAdVN0RVNsUAikeKoCXwBUSZrsySPapI4Es6JL8/b6u
mYE3FiwW7Tqj6PZbuaZpi0q+QkbXxckEzq3KpN0P/590eWF+UC940Ej2Gyi0do59
etWZTLrHPZQIIj7s1JQq3SOYG4t/78eSdOkSQKJyf4OK0juNdLsFdn3GviHc0Bc5
HE7aZAyl8RTOQcJ7m94zGqnfft9xPJxuqdypnMUjpjKcFvpkVjaO00IipA2oeO+I
fP7VHtCKuwSAtcgFoRRU4I/9/reiG4wBJg5/VooLCG00vVXmoyd9DXg9d0jPX31b
02E6ET+mnrgGLctNA5CxAJOobx8oLTT46VHuNRpEKivuOKU1gCK7JDtmBGM2Tow7
xxIvtXcmS4/bei8XqbaV2Yra1d3X+DZ1D0OrisjN5qNdyFJZ1ycUpbqS9+xb2m0m
ODSrNUNbXo0gEfR9/yKgr2gG8BqCMCYSHABoa+4Bl9Ah2B/AD2mU6k4J+G6oW4g9
EcXj85fEjwX8G7/3i3vWEsFPJE1+Y6kDkKv9Qz2S/aiVChMG+sLhs+woG+aqCz3N
ovGRZwP5EzpM5g/ZxZBXHRGjcfOqvz8u6ZnYKiLjOv8=
`pragma protect end_protected
