-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
Eacez7bCfsaEUyR6QuEJ13hvGUaUR0vB1jN+7CI+vvLr6kEK1bBFrj3/97vEjD17
BlDWfxECZ8Ea4mfT8Xc+O6uuOudxD4DqmNDVWYuWNOpkB3hXwYRh3UbnSNLxE5dB
Z2SwnirEFCzGJvwLita1hr9/BJs16zU/i4i0DHZm2JM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 8336)
`protect data_block
FjJZ7QaetYwhwNCkjuAWOeTONL52A8xefK1Xct3NCanuRHNiyWiJnToOhuz8OhHg
d6kdIBd6GhgToDgR0BbNeKYX/g5LZldER5vFRxyfv7kNnjLWg+AqH8kKyANDWnqj
/DmLz2BxqTdJijOmy1Fjl/z/h1h7i8m63dUEX91mX0SHwwfBN99+DPZ/1MLQMcR0
vcdaANdKqto4f0fgkT2HK8py/dJ7FlRjTefRCo52Vbjf5Tavog1V1VPRhHwQm0W6
Z17VLTwBGi30NQAeJbOfd3TN3L93+aloqRQ75bWb+4HBjQEO5tkfki0r2SMu1ozK
+Di53QXurVmNXR3yuq5siar20bqzb08do3pXDSzPbzuy8GwZDz3hRmo67C0kR1IZ
7J/yaGon/kZqdRVn01xA02tdW6oAviK22yRHMT96D4xnRWiefMGhytnqhYm3sigj
WNRKCzmv/jFJ/zkBvjWhAs+9s2369HdmWQfFaM3yjI2/04Wd446/QJUyWlFQ7fD/
1CX5p6aQRNqBgDUiHlWq9J9wzMYmoRT+X/5yg0SdgNuQ0aLnzUqZ2RDJkYv/3UEu
0MD6MENRIHm7bbBvqTcLkUnrMq3qiigeiFb7raUyjz4LitdQF3y/jyc40HyHRU5v
Cx5xxA2ju/+HpaGCWHC1UlG0gh4WbrFbvMT5PQhmXDycWqFiOWJFsaubl8US5kNp
KZDsLQ/NwdvfwKYt5LlCxNbsOWGRSnRR0pQxhlqYAh0jg2Hq0OM/jvya5AyI/ZaK
1yfL3WpxcOjDwxUrrCzcH8TTQSUpN/HMT/dDaLtXZRe+I7CggIXdjUzkmXsOvqTd
r0mnJ81SQlReLBslMbFWjeIkAb/YC32gCbsXP0UeTfp81so1ZlDa66X6AUo8Nro3
WBwdS/kYRU1lU/tXRaY+i6QQ8HGtvYVimBeG6zLtwD6sq0FlbKtFYjTYU0gncJNc
2pwoKd0FidoroCiuiWDcfvmI727NInIL+mwQ3nw0KBY34hxmB+xV02U3NghqgJwB
/asoucx2582M/LptFInIpSY9AomL621Rasp360xZPxmpPTt1bptFsYZ3wDZjs6Vj
OF5LnqBBzh8m6yKhlxDHQVEgqcGqpce9JinkGa4dDHpyeiM4/dwNW6y+qG4NRGxs
2H7c8TcDF/hfHuffb+sIVXXgBkzkZL+WtxJ42UwRZQ2qGu7hYuVtYIRNARgC1OgF
pY+9mgZEpEHAh+VN9Lph4YI+GfrdWDAnAT1kW94WUt4bFSVtkpeOSprgLXrcSdA2
FwH0TuQmik8NS9odnHROMHeOhHwcqPR4E00ZSoiTiyMtUiiiIDNNgU91q/1nawW5
BZZnSgoFdhTmkoq19g21WrhEdpCIp+AcyDGvOwfHiaWrPaUJQPjkzct9OccoOu89
t5ye5zahu8+3DCA1YqnnHNinI21Yn3JonVYWCp7mwAAMvlWtL1B+f2Wug2Qow5YJ
5ZqwUkNMEC4KZOShqN+SfxnNONCy3pP+mVJRAOdhFgxEpK7RIi0D4uog+XHsxEgl
WWGNBky7m5gONexdk1c4xDi7hvvF5N9WVNMqKRRll3Jzd2OQa+BQjI823dTi07X/
u1u8Yb3sz7PqhSU7H+ioFodU5KXaKxZpTMufgO2bki/vmO8iobNNUjK2fA4rX1xD
xuTbdAD7zrOPk1PcH1vlQSMDKssou4E/HM1OyUNaUJeAMvCkE1DqAbI3rKLDuqLm
WBqbXf9+veOfkvjrcr6L0gR+IP4vApkNtkKv/njm2YotcI1BBCjflTUl4fRjCxjK
+eCZWZNgo4IODbt/9OdTYAxxGedb1J5jqaRuVyHdP/AKEVNGizrCgIk0SoONFWpS
WoKYzesh+cSugjnHmwlP2Tnr8735I8zKsf2BQBylbk0jpP/sTPmkryncul6/IcFl
4JhVqDeSaBbkxEr9HCPDxikJ9xCJCugMTFOYT9y0zzXWff6VVUR6Hc41o8QS0KaV
qaudK0U55VakMG3RATZ2I+/8+VbpTrtEVKux1BtmPRnjYdAHRZwjehL8vxM/EHAL
iu0qN6JwDrNqAcrUx5cUFm7IMp6UqQ8jo68ExhiCNMCwoqDsHlDngBmCozznbi8K
e0zOeH2nIAM1r701VWiTS1pnHpLvLUWblLlpVBi2DY1vLFSynhZEVMvveujmqeXs
PqSF4dRqkztKtzlp6Ys6oqdcmhBwHx5v3CBbqsIaT/WzRheCTR7IscGsDDcufZ5O
DnxrxZ8pPfjle78Jae1d4nywOYSJN1a45kuNNkBy3s3r3MrppzEXdwNmsj8fHgDz
lG70eGwpLQMtuqK6BotwkQw6O2mg1Lfqyx7I7Wr01jqgy61EYv7bklzcFV/1Bf6t
z7qi94hKSUBvplkmlVaEzSZTXWB50aD9C83uBFEWTK9KeSb1ezuhsgbux8JzW02M
H2Jqr7qgqJ+C0yw8pqj+hulzaVwba5aIygC15JEqbMrki/qtn8+t5btQrSbmmwKv
0AHmFcpXICGBFGHNygG7/a5E1Sl/DEdLaB8SLyrM81qBDLcX7uzfVX2/Qkwkusmm
WBxi43XmkDR0fcmIueg20GU1m2e9u812+ZQ2Wi61TUjvFaUmm+k9dqT6U6lFWjFE
jLIB7LiahCNFFHnCQBNWNLVGdCBcuypTAlFJ3ZFXmdT4HJINkeHfLRJo2UcsDxuu
ChKqedaUNN+y6PJkkV99R/gUlfGPjnb/MTuAP7N62Ey6dprEUjEGHKiUu6Y/ms6c
BGqd+AOIyhiVs8ZnqvphfvEMfNSLn4OE5K1MWpdExNuOWjShLkg8+wFBlcWOC9VR
JDcg0JP+Aq3aEztrhtOOVD1C4ecDgT1xDbT7MszY/4/2ksiTEKbMy6wlZKOMCQhp
X1mC35ziD8vlgrDAjBDaflKQpgt1RxxCHIfTJVX+yaa43r9nSSw/C9AUjpFgqZtW
1yL9FM4SDY2OP5TNhzkiIs94o2tgzUOPwW77edWmmt+BhC6Yz8hcx+b4X5TmMROB
JU2Ulq8e1akEIvIssivLR8rBROO8M85g+m3PfsEaDQ3oloyz2v+D3MNtOPU4+iGH
PRkn54CklSiVqwHI7DydmEOz3rnxmip/n/qr8iRFMq1wexEjApU8hKxRDc5ibLGT
KC9aTlJQb/BC8oTpQmgtPDXq1hksNSPloneEaJ4bHbCjCiYyQ/sv2wPazDFaAyKQ
a/8YuJ0HNNP4ebSlYMh6W0gx/TVey6pYJozuyQlqbWT/9HTFfiSq9js9+ayo3NqI
RSMCorMPH/o4NOWXyV1EchVMHf2QVAruS/iR/V8ze54d6nYiJBs9biibuVWzULiE
15kIr7LDT+fGnk8IjjsOSniahAXeP9WgRHINPNVockbMMRnCRktmSH7DuXg4CrmQ
SSyIIDhGMpioA9vidsVX9sUnqGPP0yp4CxhDHVo9g7QH4+47S0agmhCmdmn41u/G
fqoptBu/0BIM4DvZP4B8mV7JmuMCfmzwUS3Eo3AxMElQDACSHfQjVHiSTJYhi+dJ
lm7TyII52HrLUrN0prhoEdBpmwPYuqRDwu4UQvCy9QQZgsk3soTa+miZ5II905vv
OBCctJA6mf46aB4Q8kX7hJUadPyTlezYntMAm0sgEAAQk8Lcccij2eN0SFGQnuZV
eqW4I14pjZsg+lzm0BxhRfeKMcof4xTboT2fm56b9p5FU7EK8FKMg9Ou/e5wPak1
ejFcCyJOIa/vUUqkelhEVfuA1969BX5AGCDxu0/4EjOvXY7tBxLrxdtUkGvQeD9i
ZOjPbUROqD0TUq4yThbQndSoiYEN7pO/24rSX78CsY1UApbWnXPMFpbplQ89snub
BllwczYTP1G6pNHJ/HUFGGZYz9lvJ+jXL8gffzLiXHZ2kVWR3K8Ut/FqegcO5CZm
6oriGFwWnErUmPD2X1SNW4XI7XS3m6pesuKkfUG0e+2683WzunB92iMhpOqsTfsm
AgJUCe5lqVDs3iKqtGjD80ArB/O07dnhLkKL6ePlcFFbdFj/sdQpDi45mbOPEPoF
sGFSQql1+MHF8E5tTFbRuYeW7dlbZACuSMaYvuY1aL8RbjlICFA4Ibh6nh+YAe+1
hkWrlY0wQrZ2egtCD/fU93VhmIGfY3RJd3pkUrH0HmesbyyAjOj1gJKvvH7iHv0K
MQFN3ECOUGQHx3muSAUuWtiokwL4f6znqOVQ3MKgCqAdBgDeR2QYqWglWiRpxsjv
zHlsaUU9hFTs7/hwnMOZrSaVF15bc3lW6u3fEdXHZZGZsP+UPN0QfKjmF5PmcsBI
H5vTt+B8kzEgnMg1Tvw/8jy/SYSzv9zEpyPfGLm+nw0CCMFSwJSif3MR6wQToniA
cfBDVgSdwzS5Gcw1n+jFE53GEd7Af4fnP50tqQMhaLE1ko4qA5t6zIX7/vwwiduB
virtsVuPqzCFWbR6UJD6dp6J4pdkqFgcWeAcetYsWxjCQyRcNXKq6ApWytMtWMUm
D19b3Zm7nhy8LbtVHHvkgMbC23cq4/yVkPOars43z4iJmBLcomnfTghONKR8Y20j
i+sKc2Z3z2helaWIQrZNvuK8WgCFTsS2cmEfw9x+BN77ubOPi5Jn9yxSWyyRUiJJ
NCJyMOGC3CYu2KgxQmzCY66Gfwezs7Z6AOzo8FfjB6mlWnqXnXCcUOzGcAmLZqwd
xJ2nyyTqHcjE51/UCwfcb8+dSvVJGhSfjS0qWzQ7JQNNlbg/t85IRLA21odWHUUS
MfvqdZciEz+e3+ufgyIV+/JC4KsByvU1d3ws4vG3hPJQeaduiWJaMfrYhDNpXV3R
wSwynBq1TqePI1gubvZpGz54MsefvWmyIQ8tt2EKyRQun1X+0ggX5lz72vEG+yYg
ECskFbzTpQjtnnme9rLdQYb/ejZgOncLZbl3voqSS/aWVfMsYScv/xMsq9RLVB4F
tivdj5K1N9wqfRYDAxxSbKimfCFpatO1xu3AdW4GNhcaJwSDUgyFq62NRiPSD5at
6eF1eS+vZ0xSqH7cbymgAW0BxAuZeT3iVa4SvUooMRqyw91EWWDuDZgquD76Oikz
kp370smH0ETPQtDSX/mvt+Fq5wagfzSb5KeGAEORxlyo3xCx9QYH1StL0NeFUn7I
wqne7BlsOViEA+Gwzd6uRJ1D7l9wsw+lECTJwXzjZtgDQe+66SXwEtERxoNUpNPi
97VYkvsBAhmrgJlNHNc32TTcAPQznZpdOffSZACtCJLKOahqMNThhG1nRLNX3muz
wP441GpSnfGcKmwiKbeSbGtXVeN2BFcqFM+rlTWA2VhxhfO978LnV/FKZ5gL8JQZ
uWp7nYklIp391x5SOrMm960+YQlPwlQXJk+qcqW4EiWJnX8ZIz02LWzCsZ78TTyD
/fXNpuwws8QbymDnU9Hv7QDgwhayoRKjW73P+DS9vdVanSQUpF5penu20xpqbg3g
hrKehmcsa46p8kHgVWVyMpxsx4t+kfdBhgno9vGP4dBF5t1xq6OeP7uJJbwE/W7L
C6vWvsFD9v8SeRJtD6l8q1GLJgeRQxYEkUdIhVeg+0DT4Qixoc/To7lkyroU+xCp
Iq4Ps+/XVmkZQ42CDRdRXfo/RLzj8P52OA2DgcLxQk7D5E85dewhrSD53Nnsp/sF
vrqcxNr3qorYa2ptTASKDRSZv0cSCr+4B1iImiWpISBMWgNBdkCjn26bNZkX/hia
1ca4v/su6eLsM8wNtKwHmw0pRuQ/hlhMMICi/eMFtxI1nqyvPBl61JFsful2iQhy
5SrtuF38uoWYxLoa4mZyggaJ4yaExcmGM69sfA5KotV//L/P+NPtofhSGKqCtTM8
+4bFZ/Oc3bJ12pwAT9zRAmytQqc1do819KIr5tWR27avBaJFLXyUHo8f5iFhyO6h
TZYXm4i9DNN+Z2w88Aa2ejIJWar+qhtX24USNt7O6rjGdB4ZBh27/5z22VYZ3grC
L6+JU4ctVKbVbc0BCHPNwVJt9a5Obz9wF7vajjINptjTPXynZiDMvI6efjXRuHLo
7vDDb4tTpHdoiPMpbg0X+pA2UjwnbVRSpo2gsWvAm+5YJ2CU0o34DxtIwfXoYYx1
UAI1dC84OOFOTBKDUzrYfn5xyREnciBFnRW2K6b3Ukg6+UapHtmBAQ0eQvO4HtYS
WcDfW0HzZER3wp4UirbHpRF+AgnhPYKnOr5m+JLlzaWdv9H/u/MbtcP0PqBlgq4g
magp5/zEkRjhgxLiqqbr6yVeHOSJMPa9fTobRfYGh7VmXvXwYERXr6s9Of6vuopX
PO9x7legfa31zeX/z/mDAxFV+bz2ikR0d0eqNYw3fAQRqZMenVxEFqTrPsQYoZgN
SpyPahKIya9i/6ETg0iQ3TX1Ciu4LcDXfQPLHEXdvfViukDOazi+2NKB81KgTbEe
TyyIWO/BvJTwMJMu+CHIPPLtZmUb/Ghxc2tck7mB9GWdKNST6VnUXabPLJkBtamU
adCJdpHXvJvxmMUTzVPFfgzWz1Y/Jc60thZNttL1IrGScvVB96rvhRYidzDZJzjM
PiPTtBZrrhwQg7dGNjHHh2jVMIFQTh7eJGOB0A13pDbHlws9LQ9e/WCAa0RF5PA6
atW1waLet9tIqpZN0S4FyNdW7CpbR4+DX+1A87oaeF8reyBLxOszovlHMP9g1Sk3
Dry2BeG8vsniYtnGIdK7LRsot3HVE30qIisujCq4qnGS3GhJqPo8HQOtpToAfW9J
FPjs4ugfN1fO1YB7TETYvNhtkHG+MB223UWTaTU6oQxYbH2+6pTDYxBxtE7IaIHo
U4MGVYyBIIZj7YIJGX9HbUkrdRVnurVsEQXNiATcQTOxZ9P/AOUARl7SWFrwn+fU
zoE5Kz6zyZpl+Am/8a40Wqqo6aLXZV6HjZzEKSZJ8XQporQljh2ZocoontRIf4f9
UPI7CUc+lm88rAIVPrnJiyIraFVx+lcIULOYBywOpNhWMQdFZpmOQFHSf9yRuyem
GBl9rsodKP3TVZ6NBh3VCpd/qaB2R40x/tWopRpmuyXvD6tahYNxjmdg1llHvxJ+
najdRXrVyD4NrRuX/wBlstLReAidsRvLnJgcbFYHJSbwbpOQ4Dixo9EqKgw8K70b
+NsmFaa3de8bI7mJXm4+tPbu+OZSnSfES3IOR1Qx5dZ+wX6RA71aGrkoIX/icoRm
Cr7wKaPgX+eNWJ5Vp999Degpds4Lv6+8Ef8s5LxU0e4TRKIId6C9RSXmlb2hcfSr
j6OlKu3epuaZTM8Vb+nl3fayVrn2/fS/jjvy/qXyrm7weD/Xspbdvglwom9Tz0yv
U7Gb47EhDxlaTfNXaHlod0vQ2AHdo0sXCOpDKiUpGV9nKGiKZchdciCu7aUObTZr
dksbW7VjRVjKIrUSzi17S0lCnfD7U3jgj7V/WYC40bfQ+M4SA9xofbByRlZ6yfGZ
0eis5T4ni2xiir0RapOMS+3Yt/i/HGptw4+Zwjq2sjdNX2srGR/dtVJmz9Fp7CHa
dnthcYkOCuiwmmYXpcSTvmw9nL2yQB0LleKzuAIK0KJMrkZqPTExMJDVkHyZxYa+
ImDbc0FP1UwWFNI2B39MS9l9c9U1LdYf4l6+lfe3CiX++Qv+Rq8oSOaeE1Bk1Yk4
Wf5iGpQBPuBu0KVGDj03qRpTlozl48fYQ2lD+WgaZSbE4DHHlxtkpSDeWyRROcbV
P2PDzZkFUK1Uv3DHHbRgD9k7cb+IUp8tNFTL/PKg1/XqpC2EaJYe3vOySU4Pun03
LRCOltvWsEhJOuE8vQvjWDOw2Xk/6WEYgCBjXYgYqfNiqzaj587x3XeEHrjsAo4l
7TFf5ACvznQCrhD4twBrp7Yk2r7p8Q4VKUjphNndJttuOeuSGKvT5rFkzahzGWJb
Tz09Vkr4Msvo67SMVKnR3XZcrJ0NRWkmeruCUOhg7FQ+Tqet1GSUa4LiGmDjKOQD
3Ud8XGpP20pBfsZENTut47wA4aRyY/Co2fnbSjE9y4xvFg8Nj8TJMIH96NN06GKO
MxAFVS1erS7fKAcRJua0prdpZjLSlVAXDGyuNQeqFx0hXHtPOhsQjIr5b1NZAbDh
x3MwzoNDdL45dgZ7NcsQE4R2GJvA5fD1WlxCfGm35uYXXjdwGBg5NlnXs1ybyC1K
ZQYW7+HLil7E69A0pXaCFbgIkNk98ASW1vo8xZKPvzJ7ZM8ra+kJ0U4poXG6koJn
s+7l9EJGRVIlt5X8ialgTQEtaiBVxuJIL+9uFzYDMSlr6xwH4F/ftqL6r5k3TefI
f73tEeKzzZTgOqH4NIDAj5PXeP2MamO61nRXm420+q8TdOTF9LECBQPnzt6EaxIQ
aMXxwx5hBksOqut8LDWMxdyMz8ej5HYcAzuzgZ/b6N2yzhKeSuBqw2xLvBiVBY9L
VRYLnbpiRcTukRV4MBq1+W0LGejDK0ZWOHJQTjhDyd8IO3dNlvNBpioScrQLu60a
y6ZB2/p+q5soTTiCP08Gl1u2OlGs1thkPUAcuMd2/uP2XzWozAcw5cSGUhCpCabj
g3JRekMpLagN/+za+4O7dbdv9g0ZGkJFm4P3iwUZkq5NnGWYevwe/kvo5x/svdiy
scOBaKLCEE49vuHBCpxPBBfUW+x13aDxDMMkVuIQVO3zB8hj9ml+JE/fjJ1So2lu
UFnjCqUZ2H8wupvDOM56h6GQP8+j60kT3deHNrtlLU8t0HWP2NuuVWH/cUhmX9Sz
A8nfiEWW188lhy/fCqg/Nc4i1CgEzdTmc2SSBUYIoVZAhCpXckeeEKJTA4uyuf4U
8RfhfRT3xkCroNZjqEY/+In7ttKpbaKJnQaZe/0MW7p08y7AMQm8E/Lh4iYm2Pvm
jxg+N3/lQVQZS7a5M9PbDeHvSBGMAEkMzU7qWtFj9jGArx7FdjOsNl4D0lu/WjCG
8ecpVjXWrH9FbzYWyr4ANJf+xbT/2Nn3SWgIRcXBoTf5Ws3WlLxQ2H7kXBdiz3y4
PME8U20ZsUlknP84KkRkTlAQhL/3rTP7s2Y57L4PQ4Eaf5AWr2vwUk8M3QsVkPEi
cTKJOq2MqVN+7aWVL3vDU3Isxc7qzzeJGVVQeoM3hdjyMW++g0Rn541ZDO4TyTWD
QdSPuJBEAfN5AxjOQ3+d+zl0kvzOIRKQjvaP7kWs6sGWWQBubcPXoorA8K+X8lwJ
rDhn2a3rtrPhsOyfTpbRFq/bM5qq5+ql/Hyx4s2lIW7mGZdR/5RcgeaJLozgMLwk
InfBdxpoPBPiDVp91sNJRa3eP2stfkAlGG5Xiun63LXoQ4SRfRVOBnsbdGPrN1mU
AcdMukXnZfGUqYecEhok+oNlbxo3GycD21NgQLziZkYg8Q5zL8OxlcvQqHIbhh1O
onn9+X4Qzg1yrvGglEOXkQ7xD0Jzr0/8Z/aTG5lqKQyHeuk4+8eRP8jf7G9QKw3W
y78K75nODzM73bOz+sDUgLoL4xaYBpdkgygdNoKyo7HrNAky4mSYBvZuyp0qPSZU
X9mWxFAamGIcrvDZmhVz6OxHGmz5NNkxlHo2PQZhh57YxzYOCf2cVggfPpknW2n1
R8+vQPSrpES0wDn/EIM3QnfvFk4GG5qgSVNB17Tt6W8cH/i33BP+aqvLNsWcVU9V
Cjlak/DdEEre9fSXbCZdjfFo01k8OW65//2Byrb3ESirmLphIluRd80E93hZxjnU
U2ggL1uMaICaLYCap2XeX1wuYJoB7dPwtPrQDXoPrMF7WPPQaNVpnX4FIF+nV1lk
YKAAV5jnOYZpgRPDQPq2YmaG8dtsTEx0d5tEIqZk3nS0xmRcCfV/OjG8ux8V4kcj
F6xVVahU6jfA+Wh3PaPScmxHMeGyOePjBqtHbWGxf5aC5KrU9dxUKR2oUTx75zVV
Xv2WlnouKBYL+0+is1iVZkHtwrRnYx/ic/Vmoc4ENiHiJonZbw/TNl17h9a5xETu
fSc8nj1GJI3VvbGXp+CXhnTL0fsrlf2+IrC8L58fBKOLBDuK6ei0cU3Pzyx1PD0s
pAQChFOS1K7q01yh2EXdTpRuguVMHZ8z7myONraHVf/xoJcI2XXcHtV0m9XDDMs3
GmeGkTOiZ35jdJjCTI6QOfpDaX4B7xXwcGaG4u8R1r5gYJtMyLmU2m2h/94FBklh
wuTLsCafeOtwds11Agy+ikXnNDBxDax4//QNlr/zOg7Z15OT1DfomBz/fhwZksJr
Cl13yngEHiyGB7Xy1ZTCI6yA6tVu7TUGJ90L+CGp9jlOWSlKrcKHGHANcH3bhKjj
A0fZTr9qJ+YSB7pXmnZPHgI9JMjD7lwFLmbA7c35FFu6qFIF4K/Ha/UkSOqtB4W5
PTBk00ZzmK+VR1ACKWJAv+85rhFJA2k1hWZjb2Sw9vbYRQmrmgpjAPqgtCgbNGyt
vr2liXKSEN/oRk/p9dghAFehXvghztGGAGYmbE7WKKQnslo8OdGN4ZHXumt/2kJk
uSBqaCosValqFqMwueL8UyQYUsZa087YxDEJeTrE0km8x0kuTv3jUp+teIrQQ6+3
0RDh/tI0dUGRdWDkDuUe816F5kInlt+I5b3mXAf9sDjy1Zw7Q/P6gmGuXPlqZlmb
Lnf58ONjyGxMIrcMJlI5btfuXJ30L7GGA2/ixJt1OJoKTMyvEU1vl19KX3bv1RIP
vAMLYz3eSJbrkqBzPZSSg4zLgnsOxIow+ZszPbtLrh1yaOoieei3x45lv+fGHiYF
bJMQllROvh1fJRh56we7xNdLMZ2rRS7om2TeudWvumKXnzaR+ubyS9OAcoE/Dpif
BG0fAbcPJEDNdSJ7srZyNwB6VEr0kCHvlKX9ccjs3nNqVEvBhxTHD9n9uetCyTDK
s8eouEqeft+fv34MAWqITBHV+cuH9+DaM1VU7J0t9IAQXo+hCXanR7FWly6Joerx
uqcSDGq6PmNsBYkdtabHQoYanx3T0MmXpIviGSNccPcw7x51VYAGyfy3SCTUtlzN
Kp5ejsHJu5UB9A6aqpXlOZzj+yW3QZs55b1T2RbhxYs4v0gL9ihpqMVziNpp/60x
xMqWYAvAJX/s6OcOQOO5+2f3p3SUxyRX9+/v2px3mg4FwyCY2xKUxLs4spfr4Whm
qf/6lB0c+qF0dMeJAMlZCOvBp8Rmv0D8F8eyPhcY4zU=
`protect end_protected
