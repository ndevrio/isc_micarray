// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
HR5F.>Q<"1O2/B)1+^OA<8_6,,%OP1QIB#@B'FG'D=M%C&]?9E)L5K@  
H$:5T,)']5R!K *'=2VY(:U0=*&=/#SE_.WGC,1>HDFFM8N]AS$QR+@  
HY>ZKXT:Q@R1?P[Y&KC4/G](GW+#P=-7T@+(5=6&YN,4(Z%))-7]=$P  
H)!O9).SY2XH/:<'[\7FV^<3Z#00+DRO[<27<CP= C"<(S+.Q7-X&0@  
H.#)B=X7JDO)#A2T0[N>=<OJ;Q7.EN?<;?OAM:>D?JEZCHQ$SF0FWW   
`pragma protect encoding=(enctype="uuencode",bytes=11200       )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@RT;,9Z:4Z!@<&8X].//H:BYE#-\XM%(F)>&BR87\_-D 
@6GVT*20,=TQFA/H[-,1"?;AD::_MP]!.LFL74.7:U-( 
@/I'^&=I'NA>*7.CO_"2P@CZCSGNMXCFC\1M/%N&D2]D 
@87/0TQ*/7W!VE4.M"!("2-[Z3-_\'7<C62TY%3"69X, 
@"A=T-<]79 !QM"+/&PA=+$T3IZI*#8=HCB//4RM2WW4 
@6J4(W%#U:J^R;C"2?WQ$7[^^)DSV ,HB9DP,@=8^!5\ 
@8@U/O^0*&28CN5Z)X2U<++M6:IN$8=V#DG.G!36#+]( 
@(-\#)\S7(A.E"E4)86J0_ J\^'*M0_PYA;WHK3.H#[L 
@DX&;J[QO*1IATF27GI(^6R]!7J3+C]9L@HV=_%6APR, 
@">%OS6KT4Z'.*?7' 3L^1\KDD/*Q7S_^C*AS=.1+02L 
@?BK&J7"%I?-U%0GB6^>D18NI$?%.C^NWBX.P1UU%WH4 
@M;8!<FIEHFDMDPKB4/).Y-I-K!UB6P9 ,D&>#M,/V_T 
@0L748;G.!U#.B>6:?-AD"23R.8=%L><%" @-8A)90T  
@5+N("&1C$5$0&CA[-GI'%(TZLNNW()J?.?S=@!;C>Q( 
@JZWXU[(.RY591-KC>+;/V=<<LN=Y13(W70J#)#ZUJN< 
@N&#8=FR1<7Q>-Z'1Y Q95L,G\B1KK<X)-H9/<G;.PZ\ 
@*JDU0@)K@<A@SYTQN?^BXBEB,8&7W__H9;_;*L$ ZY@ 
@SWSQ&"N\RV!C_]C;4)/;%]L+J<M/".[H *>+&[$B5'T 
@L^"/)J_LXZ8 @!K-!4Z(YF2W#[SAGJ!3RZ J'15 )MD 
@D3<'.C],S\(.<Q?7:V$,*KUJQS9C#@YPLPAVN%C/X70 
@=[3R0,Z&$:WD!@FFOW3++I!>1"&L\&,Z\%:2NCAHD$0 
@M&/ &+KF?RV\SKB.#S(\M7KLG<N=*2R.YC:GJ+3H@@@ 
@0Y$@UWI>"O>%$8%,1U64E%?X SII.R*/K ;X3E@H=1$ 
@(YE<[:_<0E':U/"73%ILAYVW\HXI53M1,<#(Y?KTZ$D 
@"U):M7>7L3*E\KUP7&=!BV_Q*=R%E"@X,<^#@OR:%_D 
@!X%=!.GXO$&^;SO;.HA7MXG?KS%*N 'T,)%^/U#>&"8 
@&W\*OZOM.D!$0/5FX 8S#+N<PSQN&$AM8/@!G?5F)'4 
@#3N8(J.=*MP<(+ "[DZ%E*'J6GH:\PNDF: T[U]RO*( 
@B] O;(0DDAL]&\W!)I=9'ZLS*U%C%]KZ!>PD80C3_O  
@[2BB #F/3"AR-:=51>@NIITA:28M^4.%>IPCHL&6.C  
@R/S3MV53?CTDT8,XDV$WN<S]19-4W5AFM57^E)Y:LLH 
@I,%\I 8<'#$DT.H5"<5I/1,S">AVD")J/$MT&-,Z9-8 
@W5!+#J(V?D18W4)4N*U:'="C4)5<W\+CH70?AS]MO_D 
@6TYQZ$P!"&Z=V=[S4K5(*BF[D"!CRBR-ASPE0A*U!N, 
@:9S6HJ).*$*BZ ;2?N22I;"EBR4UPBD"Q* :XZ,)[R4 
@'/KK8,DR?"FF(C^?83K-+1;_AW!%^;Q"J2';@3*#;%( 
@PJY6V(WX=4:4\GM7/-(,'J+L3E3/#YP=I-1M\+)[#^< 
@[6_)[OJ$"><P.:]H9U'YHZO,XP.Q6B\V=D 3O-2(>3$ 
@) 821ER_WWK*QNQ@3Q5[>?/0=^OYKB7?:,T#(!_U'4T 
@7]%*:#V,YHI7Z05I1-*"@'X!X2P8?"/C@X#-B_X?+$< 
@>.4>[TT3>N=#80.]"[A3$SRU;EQ>3J<K.+;]^\\ Z;T 
@("$Z;9>#:&V,7>U]\7)_L&,,[BOU?1[3,6OUG3'$VM4 
@Y S'!)*L,9L+>1H#9N#!;70@4)?@0Z5M< X[?)04Q:0 
@)&@/,T'"L/L.\K9O>(]$75?BA*+^_CS\50 54.DPA8X 
@M$ KADS1UZ6B9-E>WO6-8.AAU*J-0?,?C(!3*%Z*<JL 
@"%-HE(P>D&YP1"4M&FYY!-E!<.,,G[Z8U@AR<0Q8.;D 
@/:03=Y/3A^B[MDK1<LZ1JO<%%$I\SX5Y\;YZU'25[>, 
@S(:'0:K+PTQM*&;7MF=_1]U_;P3,1%9")*)U><];7R  
@?&RMAIZLT%<NB;)3-I4BFT&RN 5(P?32[)?D0TH"110 
@R!OY+*E%*GF2&XT/9[AYXCZ'?C@9MT3R[I981WJ14]4 
@X7BCC1>M$DT1=*3L*V(T-743=;8#@5X+,0WE\PU)%YX 
@&65ABF+4/\$E?JE"A?U01M(D"C(W^,_0R)E]L_,(6!L 
@ND:6!1/!\,> 7WG)\.67<;'5(>2K8[[-K)%J&]HK9B$ 
@#!^X)=0^<NIL;I9'2W!JF;LI"?[7YBDKBYBQ0 ,*A'P 
@:#XSUN;B$SL-<TG9YSF?$8)OM6)+";=O4E2X)"5U-:< 
@U7D--'3A.W>'U[M>D.)VHXR.F5;(E\/L<N*#F&>T/3( 
@>V^RRCQ<D$,4M=M0*_17(2J#4QCREO!.A-Q'Q [6.,P 
@"R&;QYH:"TSP*>\X;+,8>/9956+OTW)W?R4;P6%Z1$< 
@^#2[_4:+87L!/D@A/,$^*G(S_[;7J=W"9R2V7$K&-7T 
@Q,)._>AM.-_E[YG8Y<$!5C&?HONIX-ZU5O,[5\F]NGT 
@ Z*L>:*=1)>-R&F[N&.U&)NH!/[K9-6JJUQ*J!7Z6HL 
@XRK,)=&=YJV@3:U<\D-$ZWFO*3G K;1"N+XJF6(I9=  
@ZMW[@+?3:5OK@\OS1_OYH@V[G;,6A&S0J!*6+/6+(=X 
@FFRRYL$?,"0*PL_R@QBPT=!DBG(\,YXCT<$IWT4%I=8 
@UOT69E90%!66LU)YF!'/=#895>)O&=#\$9613OH7IM\ 
@#UGI4^<;>9SEB"AMD[34)%>_R_SYB+'^'F,HL.GPQY0 
@@A4%QM7LH1\+=^=BR*<4#]QY"7&P6EA+/P5G7R\RHGX 
@#M;PDD>4=T/Z@(,,&$T!76@T3_J"8#"HE7^<F]&><9D 
@Z4>#!;\GSWH,FDJ)%[F(W[T&PTX+\H2LA/RVJ0Y+#/8 
@:P5776RP4X9LZ\'<KLI@QLQKTG:<.F0D#&"7#.E]-9X 
@:K6&#))-$H4#.R959HD/#2R78=RV25;C)W"G\#Z5>4$ 
@4W+MT"4U R&E@ICI([*=0FUU6.UBP(@5O%VRBV6<[*L 
@)RI\^"<8_";U=_E=9U2-!]M J](G1 =7G:6<#U#&>WD 
@=_/W9)-S?Z<9V4_\&RC$"V4=C^P2Q A )CB\8@8EY2< 
@5F2JX'_Q5?T>#HW^Z,GX'!E&MFDQ8>HYH&N/6L6F6   
@EAA5))P(:2!%(=N*/VB$@K1UV\2<>BBNX(Q.Y1&=%N4 
@-'G(+?\<>5Y5"KA<NIKO2!-&5ZT_N9CD]RXUIN>GOK4 
@/=+=HRQ?$/&;MO5>^ \$439DY*Y@ H6-JLI2HSK60J8 
@?'B+3B8;!(J7>=5G6:IL5XQ12H [V.LE&/*?N\%D[EL 
@O:6SAP2+^.$-67F\&VF()OF=WB$?.1 5$\%DY\>\ZJ8 
@CMQ]Z'CINSU-YZ\68B3G^)./'YBF,'Z7!$02;D=" X4 
@UZVN5D;9%M:I$PFYHGL[:4D4K0OK4<7CWI2IGH5Q,8, 
@T+<D*F8K)W#<,UI,H&IT7.P2P 6DMH\(A'6F&*C=!N( 
@#%OXJ)#2?WDSK<GS;>']5"^_A+29EKY%'?';]35=K%8 
@]T_7X^023"#(PPK2Y]U>S]."^IE%8R+#]D^5(SS+-K, 
@FFO&."E)6SQ^LU^P9X8-% DU)LN_[#M/.#!G:>ZIHE( 
@U'O/N=0"Y;^[1,029YVK^C0A+&NY4 G4<KC9O9,F^A$ 
@97&G_+DD%$@0SZ1F+S>GC'/AT Y:AV'$C?%"C<!J"H@ 
@.:8W=9\3Z <7S%R<5H,71N=/UD7<AQ!&]52I^#F*0]X 
@62<#A2(FCZ[+,I*!XJXV-,!2)8BBXE"9+WB>P(:=1,  
@!IL!2+_B->'>A.SQZ#GUV KG(C\(^\,WGXBHPZ3)S!$ 
@\3DTDV5IF55:VWGID[,T#@V2]!CKDW>^HPY#(WIFL3L 
@]8FEZT7T,@@QR)_R@<)N:_!I/<+/TP&/&"/$Z<E<A.8 
@X3Q:&\]!KYDY2W-^@="Y8G7>>\;-F_8-+$MP\+:R4;L 
@2)NDHK-U6WQ.%YRN567@YXQM"5FJ['*+/P1M!WQXJ+\ 
@]T?8$$%N6AJA(*/XG):(<@=@6^]W__2+!6R)*$0YLJ< 
@N+.U]^=D+P)$RS_&#:&$C_50I#A U+17]IL0(AV$^2, 
@X_:E!]?IXZPZ[C[>6FG6E505U'QI$0\PZ3M+;\N^>-< 
@LPPM%I6C4LYV\HVFBMGK@45/1]#N$GK JKGCC0EK_K  
@VN-M8[:7UPR6.*,$>[YE;7CY=[NG,F@27QF((EX5AR( 
@"N "S5@K*IE/^D2KO(P"C3WFR0FR3R-BF544((Y3R9  
@B^H[0)-^S4?& P[I4!NPN*!U>,S@6%6JA!YN>,6X,&X 
@&9R'EYVX#6'BH"3_S"9Q3L%W9V3L5(/I(!:-9 0C'LD 
@&8?$VPF)M@5<HJG%[5Z@G>&GV\&X4YKCE^LO:HCUYLD 
@C7?]$/3]YGD06.K,F]?3>C% GXA)1O-0V8+2U.%0$%D 
@!2KD':J&^^4R[FHQH''FL9=#?=V,Z(^^(NY,3PQ,%Y< 
@'_A:QXQKHB%)5MD"O:+#16$!YE#*;/7LSWA9UV(4:?0 
@D],/(05V#N:H$6$4H7O- TIM5NBYHU.]AI8/QF2M .  
@J_T(/;9 O*[N(8B/+8KP<Z8RB4,X8,]KAS-'6,R5BDL 
@#^&HD]',JQP:3-V%M;W+)=%&:#PC3TAQ8A_M%N;"RUH 
@E:?B>L+][M[!#4ZF:AIZ@Q)%H*P9,;H9!D2'P6AUD_H 
@87PH2I0//PZH(6)R5SYZHI'\]ZLP3.?9(T=<VJ:8N&P 
@'\I,/[7X'LT"*A['3>_ F0C5"&WLC4SO&OXHODI'=4T 
@/"HIBMI0_C-,]H=EZ/TKL"QC,VCTYVR\2<U;.&,>F+4 
@JSV)14E:6(QP-KZ3II"Z ;DUGL%4M()9 ]VYM]K^P[H 
@U>!; @VI6JY0$)O6?.,\HJA-NT*5$FJ__1]SVI[ 7/D 
@WS5[T9A@/? CYQH94G"'Z!JWR707W_RU!.S=*"0YFHT 
@ ]<:T]OUAH<$*@NJ>'QQ)IPF(T(8RT4XZ4<EV--S.CP 
@B R G!4YTWC%>9#TO7#9-BX.7;8H%84P#.$J /6I/^H 
@R5,<DTA:3>(;C.\Q">.0SK3C>2.W$S8\F"7R3)YZ\8D 
@K8A+P\]1QO >5<-;3KOE^BORM%C2J10@)L*:OSB(B]$ 
@EG#$VGO/+YC32-W+0OTC )']]+2@;#.YJ?TZY62)I)H 
@?Q")0"X*#,#67T'_<ZC"'_82>._ BAYT[.D1AZ;-Q\L 
@CV.0H4K@$@UO^17-@!6:K,KUZA.XX+@-J&SKE+;._I, 
@71@E]0<NH.0\OU:[ZO/J2:OJ-78\@58F8VZIN*B:B>\ 
@BD/\F<G&ZQMQ^F^['VGJ\A!D(2"X598AT-(19V4IC?< 
@)*C&Y]U"Z./I@$]ISX!A1^1$(D\*2,A22;:#G_S/N8D 
@MV4G%OECDJDO1B[,J+Z2&1(Y-6IAYX6_52?9'NF_+$  
@\]9W[UWIWHM9$I*71[I @N?O<5DY4_N3NO8D:PR0!#4 
@E66B#T=9Y2=(DB7FRAI?%/6WP^SCVY(WSZR47744.]@ 
@; ZC+[VX*6V$ZC1ZA;P_E8YQ 4S;?9>'_X#5I3-4VR, 
@\,AS-O8@;E>TR6(@2H+HRE-PBS44GPUSZ!(A;X;55E\ 
@9&>F=E(IZ=A92!T-Y\"5=^WDVVAD<Y?H():HF(/"LC0 
@B$C!'AF?7H:K,%@EVT+ _Y2W_>_3["%A__^#$NS$A/L 
@"=FR^/2#]A+[>_+#BU@3DT@%A"_F,LK8QRG&,1,S+=D 
@PE5@L(AER^ACG&^'CSQKY$?18K@I$+%6SVYV# "B;#8 
@9>#8RX^(MBB4<M6XP[/22U=9A5)?0H;HC<)5<.&3C'H 
@.4E.L[+"3()#QH?D<:9@7YC%VS(X>*]L[HE?&14.61, 
@"-$ 9*X.UU,0U@J[IED/8-#1,J#1K2^H\$8O>.E"B>L 
@QE [SA+&3KZ]3$"#?YSPQVJ9(R*IM^-MCNSN=)3 P]$ 
@]WQQV__:5<#6W O=VMX87@:H3WZHT[D=#='1'),PVC8 
@_:1T![$S;Q:97TGK+]*N6G2]^=EK$[(JS,<-EE:<S+4 
@G!AG3ZF$K>GNX95@"ZQNZ:?(#]UB5&R)Q$NB,]AC"!P 
@Z-K(:+6O[X!N/"Z(."MW-]_,;O$X/25<%],OZJ1=<:  
@L4J+JGN5Z[")_3RB9".5PWJB2*K;B<A0C#9D=TUOP;@ 
@R;N\RU*'.$&Z 20$F,^=(0O<U2Q<T.%0/F:8$8=BP?< 
@G2;;S(&Q_TAJ!."DOXF56D3PJ>ZO%V']=DP 'P4)NOP 
@FT052X'E+SYDAN=D3( 5KI)K;96K$*ZLP)@<KC( 1N$ 
@L8@DA>-$Z.UD+H=.SG)[%"H\,&A^,G1P+9!,2<-C>+X 
@WY4G8?U8N6X*AXFOU&=2#?*&AY0)82_6TU>V:*Z7H(4 
@P[0C^%@#39_>\#&0)J"8<I?Q2>(:TY_T?V>"(VEFYL( 
@DU;"[K4O:%%CU)#NF> ]P_:*&^3OB!$%_ZM4R9)[&2H 
@1"0DJ$(. ANAMNH5,?8PF 0 K[7<U&1JW$'CW&3;E7  
@S'29P+FP$$2,VO0=:-+1^A[S;DPHBIQO&BZBNXKZH]( 
@0*L!+RL6 )NC7!J%XQ>&(!8_L!P #T^3[ C:>@U"$XX 
@ZRNQ=67D7S\_=:3U0H/FUO"ULQ 6\R*I'?]^_79TE(  
@=&YQ9EZOIM$P1$)G4#/H8WPPG#JGO61JQF;,MQEE_ND 
@;9L6$*G4_G&"F4X T'"K]!BK*40K,E$'G>D7A?YS\]H 
@TR@4B)@9L-JL](>%3G#J$FSYNX%6$S.MRAJJ"</Y3;X 
@\GR$XZ5G*9XZ.B0I=E"WR::PN7@\ M"7](-03!T#4!H 
@J_AE6T,W]GRA22\>R29G%ZZ2U7RCMVE@K[2: L3#X'0 
@15W(ULX69 6C:.BMG&P*G1CY,=(S9MI4];%LI:8]]C4 
@W\NN0;TP@4N+^0DV9^\4+L4.>9C9!)/C70!B.;(WJ]L 
@4@>IYQ<XQ!Q*PBQLE),CIBT6%<T5)KI)R6L3_+0N/?4 
@[]X335/ *6G:ONF7>1>8I:,'M0<X+^U50_6:#^KV<_< 
@,D2HMM6/GB46,3MEMWR?E1PR0MM'OY#,::#DP 9#)L8 
@$935=%0]3KGI&L3%+6HFSVQ@;;^9=+Z$*:,MAO@0,XL 
@ZKH7SL/:;=!10;:"++OD5MA1J:/F89@ "*9_U;QT-UX 
@75@V.=XN?3CD1C=8$=TSHNIU-7%_2Z:EN&CS'K?YQQX 
@-T0C4[EWR-E&%7]-^SZ.4JS<1:&RL:(3L3><"N&4&3( 
@H&DY0I[B;5*H9MY'Z8$&WU_?C+EAJLEK IKRR+VB; , 
@#.%"$NF(0P=&1B!GLDC7WY$IYS![L1ONYAE.>&_X>XP 
@A(Z&-*/@)6>M9W:L2T\W%"XX@L.WE=,")5^SF5!V;K\ 
@ B?>3SC_KV:53@N(<E:]I]'!ZQ$'?Y4P)E>[!']OD\P 
@GC3=0T(/(1PATNL%CWHU@S0<#DWDXI^L& Q+G>U"7PH 
@XT>F6LB\N1W&L>N\ YST1/(7AT=YRA?:B5=OJ%AXO"$ 
@.]&'O]W8F5:MZH=/@"ERQZ82=$?1]WWI76LF:WDB$&8 
@F"!^1J0#VZ4N@:<B^OBKQD4J%$1UW.&2$5/]MXE=B\8 
@H[8B 8C(8*(-B1[(\%8\OXNO@H4D$Q@Q_FE@;=&MQ^$ 
@.N!,=]@6!&I=-<H @*J\\C/L=O,E[]]).U*:+=_=,7@ 
@R!#=+,<N9RABIQ/S].\^H%ELVDN*O6$8NH-SR*LS_LX 
@$7=JJO;3#8 !I?2-+^Z">M0,&<<9SAN^\.\//0,KT50 
@_V^-E&CN?;LZMWY0_"2NPI!Q0':)AZP)P+^(8E\0>/< 
@EGA!TEJJ*D7DM%.51^_+1&MO<(.Z\P-G*;];B!+&!Y4 
@R-4'Y8!<&&701U0A()*PA(WZ<)9[2B*/Y^O7%>A[7 \ 
@8TSX>.ZL!L*9:M& 9_8G%F"@JS$GD_FMY/\,U]NCM)L 
@H2*9!N%+'7^@M]:A7="O.$E1).'?'DTAJ?G'.'&<I6$ 
@K[QJ\H^P%BR4LX=.72\H95O=0U-^:B*W0-8IX=,R@4, 
@S24;=CXP6V>2U;?_QR<6:X>3PH(64/&V4QY?)=L*.;D 
@*7T-8]O+C48QH6+/(EB5[-?X!6]N$39MA:HA9#J/+[\ 
@Q/I#+&6R)H_5YRK?WY0T<Y1LL)Q_?YZ)=B3#1V=7H\@ 
@$*<7QR<5H-![MT*BT(MJY,5>H06GS_+ E67ZZ+8RWJ, 
@?4$^UR'J&\X\<"- JR_:Q[K/W#XCFL3(3%]?J/,[@_@ 
@@#)KJ[D\- HJJ%D!^B<"H$'&.CXM:34RV-4'+#B7(*( 
@<9KM03!H ^1IJ+Z7ORFP+PNS]+B_BB?7NGO)I1D?>.P 
@%B%"@6TP?TYW3UM,X&/;AK_D[F29&]O4ZFEOBGU%C.L 
@3Q9-041?B(\V(^'CM<@N)2$%RRI@0M!!)7JBA@D<<6  
@/@V/L(4O%-!=6I4UH/A%.%[#2)2_X!6T.9@ER<FWO/0 
@ Y"](SQ[!JI<"&H!ALT\NYJVMO)6>8)A'49CIH0PV2$ 
@-Q2*L;!;UI37Z2D=G)QS6@<8X5"K'GB:@MT'^[':EKD 
@RTN>REHBAPYJ1]W.;)3BUD)D,'?L!RW))6?07C3429$ 
@!G3:NQ[D'=QQ<V#H45)SMCK3['(/SZ(-2&I$5!=F?.  
@62X#9]3+(?[!^>.:J$V?42SZZ[]?TA(%EF7('11HB9, 
@W(*F(KW1(GOQ1<^?^,G>PEI<CH:A@4+.7 G1"\7A?V( 
@_O:D<M2KSN(.:97;BT\U,\4$63#]T%CZW(&Y?RGO4GD 
@,GM#3DOVG 0C_K\T*F0Z!:-NHT5.AT^#L+0\;\L"'ED 
@'MKV45,\2"BF0#>DP4>>G]7("EQ5[MFA%&?XZB3YD:, 
@ZI3D?]C8:8X2UG%/>I@1U\;F609KR,5,'*2XH"/@&B@ 
@$![@[1NM&GU**?+82F)CG)'M)2"F;)7(VB9;[2(6#;P 
@>FF4FIR7/&9LTN>J@VA&[OY"'N",Q\4H%K5:E91I=O4 
@T5OC7CH^*S9G<+N:]MHEVX9[NH#A& QJSDU1I.@M-@\ 
@#B69T]6 /GIQCB48!H41J X(5VWY*$6Q%/Z7U3' WM\ 
@@V/$F:FDW,>_X#[,V%J>?R3S8BM,Y"DFE0WZB"<>SLL 
@;C,;/*HQK##%4X\-$#AG1 92?.-:.^8<RJ&!6H,YXB\ 
@&'5<A.JU>R7.FK^3_)[W(4S($_B;\>Y*6PW^ST?R/S\ 
@[^9:?+?Q;/?=^-.'VMFJZ8G(=O],WO_C#*G'TZ52A80 
@OHV<^)LMD/F3_CL5=K3?5O5WV1*D,]B18U,%XS[)>K( 
@Z[3.[9T=Q]1.%"#K8:=14!2YXW $C-$']U+(RLL=Q+D 
@PP8(_93%IL]B8Z]JK-6FR7&J%6*^?K$AS*G</6.UY^8 
@O\4U&DSX>XMV;RQ(JGDD4&<G3W#EUG,/]SG9AF/7^[D 
@%< LC;L^#\N5?JURR=>_NF=F8W+X/D&26K8<LZ(-0%0 
@6(M[K,F<H/ZP/B;@GRKCS Q-Y<B 2U6#\AR,X D"FH8 
@,O1[<-MRZMP*''%'3*G9?;G**2GT)RH'RB "^$S5A(8 
@PE6X?>U/$$AD>\(@H'B\AL[4T9_HN,ZX':2WJ+5<Z>L 
@>H&7,L>$R_RJ5X>IQA&%)9=&Z)#0\C%\?T*=&(>^D>  
@D$D[+IPL0 3^AK&G@<. -BDR<QCA0Y*5+"UYR>N"6<< 
@6]MFMVX9CHVTF?K:(!>G[N= =^<XO;7& SNI(3?XDY8 
@[KX\65#>.)DV'>@*TV!!H"^4 VI'M\!<?3=2I XB-.D 
@AH?1$TA-WGS44P=I0$Z;2.)RCYT(>%!IMHW''<2YQ#\ 
@2@W6LG('#1(E.AZ1I<B/Z+3 NM0RC4$YTG1:P;>?,IL 
@_Q$>;ZS%1:"^OBE6U<!GJ!?H+_%1*YH.\R/G%FNZ%9$ 
@/2_-WMK 3T9J7AX?GU6MPCK#4;(!7J6I^?N'.2HV34@ 
@\]IE 62-:EXV+#_[:3&2OX9BI8)XN)VH9Q;F2"]414@ 
@ Y"Y9Y0H8G!H<%E\#VT<0C>K\RZ/Y$0CEM]>=PKEB<@ 
@(]$.=59X+#.22_*CT@3#!'_?2L'.VF]$/=R5XJ,-28, 
@&XP2\>0RDM,.>?$?KZ$CY_:5$CGB(P&HCRM4NGI:E3X 
@&E7"D^O.3!.C;^SP$61VSM;G-'LJ%*PDUH+]K,&D0!P 
@] %B6JY566AS#NF%(%N].(,4*A/:0F; 8BJ:PD VV7H 
@S0(QC PN<38^"Q0(M8?H;"L#ON[IWE,2Q&HQP&I(N,T 
@BL4]-.R<5E&0O<CGMM8E9O4WM7GUFJ2?1$5[X9^$]A< 
@_D2T'R6&>??"KDAV.]%UN=G?!=H'* OT9$&/4]TEF20 
@J%-LIF+>F0N'*>&2S>1VG!T%C* Z)0QL=S8ZF-$^K_T 
@"-QRSZJ5ME@S%+;#VM^5RG8G.<?GWI?<-,SK T)FUR( 
@S;]:HQTZ#3-$,V T46LQ,.FPF_'\Z=/XX"U]6E>$4.$ 
@Q/L;S;R9-X'LOL20I@W=AYUU]Y#D*8%OY0+F5+>]53L 
@9\A380)6:A56E8D,_8^;[.<>W^I=<!S#]_@PZ4LVG3L 
@_9=+[I+TDPIG_KUIL8=G7>C'XII6*&IZX$0LK0]'^B< 
@[=P+3C-\:Q3_2Y/GMUW1A:M]SA?VG;'[IC 1[9; )Y, 
@S-F@.KS#YTW<3$6TG ))!R&PHK7-W!LFYW]NHQ% CA< 
@0SGKZEI^M1+P_OE>_9_G@L]X .9EG'8[H]/ZVG<#2"$ 
@!ZE(8B[I$;.Q[6H$QNI;^_U* '1E^Y"T\%\'KC&.7=T 
@HCI*5'_JD=2<L.:!H9VU[?^-EDRB3)557B+DC_CL'4\ 
@/KA!C_YY,Y&>)9]M4O;&3I+M1_7R_V-3E-F[DO[I6*, 
@ \#Y\P#5V+GMGM4[Z[5?;="UHS.H9!'5C^HL25;5* X 
@1]>'[=!%,^:#=6$_Z!=)>LMPU(\C"U944^\5!P9YLY$ 
@,'$P,VL&S/!5P:"):WY)B6> BAHC04?=<_^K,9SPE=\ 
@6/LY91-,^\(L+IWGZ[;.WY?Z-0ADNQ:(H?7(;V"I];D 
@!^CC"075JF=1A\+P]-Q,C44X'XA'ZN3N/EVE]/]W1/( 
@*8LE@9/KEV]Z<3+TR=US01$N?:?*'(*R\#F,@VK&9N4 
@&[D&E:8Y5&_1WWPIR,D3-1SZ\-]C]OM6\"9&I1$NR?8 
@350NU9E0#3OW^6?&L#E\D;))_P:W@*EL.:BY2RI ]Y( 
@8'U /N6"+:4Z5BE/,CYDB75 _R.[FC$"RKA\8VGM(]( 
@AGW)R!R?2+ZU\V905YY8D'-UAK&JYV_#P_M EO';>>\ 
@OO0HYQ(=WNA=3F'/F*,V*%<:$S>)JO'Q:T&8])G[L(@ 
@)F;PQ&4R[?*H06P$2M4KS>_T38"MW@^3S>UKYN.:;I0 
@NN^3KO^N1#=D#GZ@T?J/Q?)'"=!:SAR2"%M7!!EFQWH 
@KG;YA QM1JRV>2OOS=X=QFC\+VC X!H3D^I*G?-#;:@ 
@ECX3.JD*4P",KIC8>E!R&BM+9\<CH""Q^.N?=S*MY!H 
@I_>OEN_MLE^?S&AEM4SNZ\$]#2H*'+$\"26+P5U'W:\ 
@WKQW2) "'MV4CK,,(P'(1'/$Q!&4ED%S+'+9C+2"=V< 
@0_YK/^0L71 A"<0%@]2%!E#DW#A6VQ(@$X9=L!F-2+4 
@</%YAPD3T4P_XH*7K!/'/?@-1@FS+-A:(:(GU3EIG#, 
@!SW&DLH^*>R=+.K5_<@P@'""4%!FGOG1[8Q9C(Z+TDT 
@69&=C:E\#??(H6\[;!91:YK4:N:'X^/'LK+^D?+U,+  
@L-0Z&(U'$$\UP([!>^D;SUW8"WXT"P_]JE]SS3B@1D0 
@*9( T0B=(.@/_YI\11WWMD-# 44"T 4-)1S28 5SV>8 
@L'9\PX](92R,@BB1?H.(2@#8TW3.2/9,E%!FT\"(X,, 
@._3#9KO:ZC=_4H5<Q)EYF2JAF9%$:MH[/&7_%#7SGB( 
@ 5]&XDA3S@_FPN'7,6TF>TK=YV7Q5Y,K9LQ'_@-RPZL 
@+F!V#F4DV"#>+D3*Q;9JE5 XUTY^O6TIEU@HZU"\^,( 
@K.<JX5P&,C$)I?NXRQBAT5^2P4/*%8.RO,3AZ2!O "( 
@H[NWC*0[C*GPF16#6N"[\2!X#J'B,55;]#@,"!58=H( 
@6;/4IU2\KI#,9858LVC_K(FJP#3V@[_@L-(OMB4:!W$ 
@E;>]P&ZT:E "D\:!L$E-S!T23YP,9+!3%#-35-R,R2H 
@UP06G8N><=0O<42ZVS8N,9ISA&&O<QQH'!A*0.%X,.T 
@._3HT?K&8NED@[EI&@(:+7GF%F6I7<9U>XGE;W:2M>P 
@0=N\1,/_%3\H:!G@C_(% 6=01-B=O0Y%AA)&:E$B[[L 
@=0O2"@$3_6MP?QXX(LG":.AD1[*0@4+&5L/@?"KMI+, 
@J+!\^!*5RX.; I?]ZCZ#UJJ(++Y$(H2]B K#UH<09RT 
@ZR-?1T^6SK7>5#8K)_,-FO@$]A0KBHL;'7^'=[.C'/$ 
@DTI#"-2ZX/1PX)EK4V=S8D-CHP/?4@#D5'4!?*96UV( 
@/"<D^1 )D@6=_8EHVAWFAX>71\FU&!,WS6#K/FOX%T$ 
@!+T-G_>.>K8-C2!7TYEEIFG7Y(]9V@I9,< 5:;VZ:U\ 
@>C0/==GD 64M) -3NP%^4 ,;X[;O%1"'\KC1Y),'&!\ 
@;$B&_.LP..'EQ/D=H=@Q2F)@MM(SZ8N46$. Q6(I920 
@:M8)J+ 16/_7=W&^6&ETD Q5^10O%]9'%(ZM[++2#2P 
@/1ZNC1;KM:';WS9(EC ]B]C_[,[1,>@9X<$W%2SZM(0 
@&-Q4X[U3Y 4VP;S2#I4+,VU'TJ/*;?D!:6K)4>1B/$, 
@0YQ?Q-A(W*4BC<D>NQML/$89SWXY4B1;<?.:5&:B=OL 
@>(MDYKY YK,%"30@&J])/<HCU?]*5*%+'I_L+P;1&_T 
@[?[LM]!B<8 U$3++9<$^DJ XVO.LB+ 6?BNZLVYMJJ( 
@@")MLR8R=P7I*/8//30^62=_6*M-,* ?%CB93J'=00X 
@X_T265"ZZ^R3/WVO2^6F16Z^^="5AMW8\PZNU6.OW3T 
@3S0O28E,2SSR^YJ]B*Y[?]]>M9DD1IFJ;SRO1L2S9#P 
@;<\A=+O+O=>XBU=#:W_3<K(M2IZ:3DYY8R9PW;VH\*L 
@ZV(>*'H00LX3#@D6%^G6G?WS2X6;X)BOO6#_7O#RETX 
@WE__W,'FB9J=-CF_1)%6U\?7_,@I5W8/)X;8_(3/PK, 
@I YQ"F/+'D<OJACLNSJ;=:+/2OB/J]NP6BO94SMR!,4 
@:J'I/=K$5*YI-C5V@#;X?A?"*<CGF,#L&TJ#N==*,GP 
@T'!0[\W5W;(KJ (]6R[B'O9(T_QO^@E%WP8E-FH>?KL 
@$_=*PF;.;M@X$@Z##LM8VIQI+FECH?5U>-#P/%J''-D 
@HV@<!29YF8B$R;1X/G-^G#%\<\.QOZU OE5X( * ]>P 
@17R)4]!&6^<$5]&S14W6X[?R=(D"J(P3HYN1_Z31504 
@D.L,$7DSN6C@#3?\OZD95VM"I-S?QND7LAG(CD<F.FT 
@82;2WF1MJX"]9/0<?]6B=:J%>Q4W.7';06(DK=(@"NL 
@'I=%I46,ZQL>D1;A>$"EN457,4Z#+/);,<VZ^5.H 9$ 
@0J']5/2EA"=,REI7[=D!?RP?3X=&Y:L:,/A5KCLTD-D 
@ *B@,H=9BR6L%CMIW[D_823UAHP8.:BS]4\*_IGNO<H 
@>68N)HHP44MD%&9O[6148$M\R+BK#<3T2ZT9*L\&^MX 
@ //S !Z[!%U_@3>D:TO,)1_#<N\B=5>1^\*K1QU=VMD 
@JDN,RW$69EIV6J;>V #M&C.7&I[$O73BWITOV<TZ(V8 
@8IQ8Q_I17"E.5]B]ZH%ZMD^B5.*!?4[:N,,TZ\]#L0\ 
@CBH/O=*HH%FI#(-JRI@@?# SYX5-Z74;[/H<U(:L:&$ 
@8QM;=&I3-7]J;5?[T4##4^&P="_<(/Y;NI*T50[IN\L 
@T&_:(0@ELA0I@])5H=D+/1?703]R:UV< :%.D-0CX_8 
@+:4C(HG1]<$BL#-?)S&GYTJ JA[\%57YKA7!X%S$(BT 
@5F"Z"FOR)RPQYL!;NWPKZ#NKP6AE>7=FG^LF"#*+MCP 
@\PU8V#SOVGW/D6P/RZ'MH?Q*]O*.":$G@1LHTL-("8P 
@/3J=NC!)</V=B[E&%**55!*<8S94X;W"A$^4I8YIMV8 
@+_-:2,W44[\Z/38E9 [%2Z_1/R^9KQ^QG,N+"Y"7'#$ 
@"K)S5$92C:I]@Y9B]>I:K";\D;S>)0F??6: (WO\"XP 
@S_4UI F?7,]K.41X-GV;RMT.CB_H]L!+'6"_K I#UGH 
@PLF 3\HEL51X*'0UJ-T03.$/HE5D]SC9-I/C-"$Q\D4 
@+O2@8L1U,9SOX*R*_J\U1*8>?L\'74* J<@"*;P;FP, 
@NP[ 9&_O\'JC1+_GC[@69VYAE&]52 (6G2;B /T>$&8 
@=&A=M.Y->?CD*'O*!NT=,Y#E_49O;)PC=Z!1UO5G>;T 
@;JZPSP3LM]T<V$!!I[5*Z3THD(*3]"Y=6!I=+A=4FGX 
@$H8_XY3\H&4H[3" #\KJ%F_SH2ADC=\FI&0BBGD>%E4 
@;V5B^M'\ZCF+J LOTYJY*YN9U"*8>J(IO/C\T33CC9( 
@3B3&5;93T%?:[=F2%&6D /S?@TDH=^<"XN:I0:-8?]@ 
@G<D.2Q,('ERN8#O$O)9E#K7IFDO<$N: .A 8?>5Q,I( 
@4IC,-^,A,#>$'30+752_F<S@N2FU44K,\"WR4,;PV7D 
@;QD!>#+3$6)3OZX?J4NW2H!C>(K[+;M"&QOEU0 &;DL 
@)LD,=S<K%\8*0 VQQDE6RY4]59+VGJ)UFDK/\"Q%VOL 
@3K2F5QP>@6DS:9,\=.^CE<3,3>^)U*$X<,TG->JFLJD 
@S)?SX(XW6K6NM6B:H(R3C^QUL^]U-P\L9 O?DEA-(U4 
@QC6,$9J]==8R89R<=F:!IB6WJWL5[HN%R@\4K=? [+D 
@1RC',,8JN%4!GSGWGOP;D4#;R:\;'*.8WN^'2L3NL\D 
@^=:SW!:^IK9ZKU8])!U.]BXVT<<:U.\<VO+.5"\Q9*H 
02EN Z]760L)X)R;[[JV_Y0  
08 ,X07$7X00,P$7L',9W(   
`pragma protect end_protected
