// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
DHyh+Pc+zA+19cO0FTs9mS01tWmFVHQEHjCNRfgsgdjuvFPwavJg8KYu+u8CCG4SgM4LG8XaYJwh
KShfCRjXbUclvwrGhOUBAlXqHh8FAx60teman4Upq+RoPgOlkp/0HWiUpubKWzJknDu7l4sNBYJi
gqVdt52x6QjE8x98mW4SdWD0UpVIoZbbOGpib6Kjlphbrt57Y7leyNZV+7TesUmhsC0Giy06mdXh
GEwpE6E6eWV1x0axqgh2zgWr5BmgVAfD8xxTK9wCUCwgnUZ0nyeBhzJ+G64kXgtQdjPkqmJR7jWg
KbmJAEgqk0q/Jyt6/jV3UvDBETE4Fl0OyL9b+w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 23696)
UQoG+9EPtZpYm4lvK/1BOLPb7mzvedMyrJ9YVpjvyhOc8oyo5ou7Wz9g1NS/5LLWG1g5gMERY3i2
tILEbZVueX/GZV/1c9IFRy8bh1SKDbLq4vhtBhgcMt2Od/90C7KBonj+HqJOoJu2Cq9bGatKW1/2
EEa3caemf2O4OkHrcVsSOMakoOZN9N0RfcX0Qdkb8koz1+S1mfYvHtrWn2+HoIk9MLTRlbxT8OP6
MCNrwt3tyBN16KqT6ZiYhgd6bDumOz94uE6yMru4+DiwFhzt/z/ywh2Q20sG1suKXyHVCj8fVf+c
mWY3uZWEzLjTPQLKKdMwq982li/OzXTLvtD+Gw44vH4pTZWc0SGwvyHcY2mvGceLR7XsSWg4fnnE
bHfCAt9/H6T7qy35WVm0z1lalR8tfZYUMd3enMQVnEayxZkg6f3wJtD9SjBQFuU0D/kcbdewUZbR
b9mQ7WAXZoXRURpCh34SgWrFsVNS6ko05rdQFM+cgChQRGgoT1Xd7J8w9ayhL7tQY/dcOzCpuc8r
aV9GHdUg0uW+piub3VQoujAAVDPjd1way+sH+kaDSxB1aN77D3tZ8hT11hkgKVOqzHf5TaFAn4zS
SX44YMDIiyoPL7SoVP3jj8jmJBZpR412PQPS286Rimamwe7fBUsov2dCwg/Ib9KRaBzTSd6kIU84
PwgT1x0wa2Mx/Bxy/C+nuBBkTjs+hJnXxIscjf3buR+OmJMZJemNTM422MTW6Hxu+yUVRNkYdpBq
4uWadeMkTP4xhzhiGqP5wSWnIJjysR4xxWiQ5I8uk1+I9g+L+bw7PM9oMVAMfdSfeP3HwKsbWdyw
I7mVLUkl/gf62FK0Tt5Y14BpOkZhIsrl7fmHAwU9v3MZ4uuaSac+c3rx3GIlIm9ZZkqt83HldPPh
OiOY9PR8zg+xlfaoGugmNhtM5dNagNsfjYJnoMjNCxldx2YUG5EHHYL/Ma76CpuEa2O8Qb+h+96D
TEOStPDMkOz0dMoCsGu8fQQSGtQTfs5JdsOQ271cICnzOB3CCMQhlnKeBVkjXnk+Q3+6P5hLaaF9
mk8bjCgtD/GigpFG902C2qVZXsAdkjEctEtMXsHtj2e79RBrRn6kFFtThyaC5hkMEPVnos1gBbzM
OpGq8TIPGbzeq9xhWqJqp48gf4oL/EbH0Um+59SodP5HAZuJH19t2ntQkKbH5H1RUAYylGLiW56S
PmhhYdmBnhsqZzHx5+hluqsUqPtyq0Wgxw2gGQiFenmDQnX585iFiktSch6oduyPBmQUgDjOOjV4
BIlp0F9zeO2P3vLSYrmoC1UUaCxRXUczwuM/CAwmssUhQraa8GQ2KJ0t60pbbyAiSr+zohlCWTBD
sryt0UNduVimCZ0uppA8lu+rPTZq4jxEm0jkCP+LJr6pK3ZJdyTslc8rm7SaYl/Wi5a32V547q9o
5Dc0UnoA7g9/fsE7W+QDMMMRiP/FizZXIGcI+ii/pOBmeXE1hrL94LWGebuOfbR1GgHGEMHbWWZ6
wac/i2hsShaxEE3CsjogaS4FwzSsohM/TSdWOO5rAJBgi3zJHxE+FVkQqMdduPQpK9nteewDbrqR
adogYPSV1VYJ76MfnQsrRE8D6xOFGu5R3kbzBscDUS1pXbrC3aDelHUVaC/2yQlQy9a9VF+nUKeB
u6sxPeo4A4VOGpSnOQXPlAMq1ESuRdt3YTqCy6/pE4AAN6wop+Sbsbx4BsiW1g9q8bPlp9ZNwH5O
MI3UgettiKbrMQ9vdBNRhOFysWSRxTLZpoqjX2w2+QE4fRqYYeQAnLX0GAt35uj/idz5bnDW0/pY
H4soxG0b8LAyZCSj2sKaT1Pt/ANXWHJt5N3fEFO/6c2hVGLw0L5tKb1RSrNxN5Z38ID69CWZ0Thy
qT4+mDfTAiyK0a7ed0/DaEbxn5aTVGIdIs5Yt/IHb8ZGFG+/UARqpLgqF7lYe/dFGep64R1cgJ/T
8017/B2iUCkUk76EIh7SNsczXldf1GISYAx+laCYqXL1BpmIjjvt8SE1dBv7YOIhufcZ2R4LRZzI
TiOy2s7l5vIEa66jV5g2cJIQUIh9sg8LTNYC4hFw0W15jSbVBE5sBZJG/uwcpZ/lkiW8CxEpG7M6
EoNWoDkSyzUuSy6xAy+Wg1ctPBCAB4Lr/Xm6wupeGkAav1mehGy1vJHlWfm+gwuFzx2YC2TuazKc
M8urE7F8jpbgm395cvIwQ2Vfb0hSp4BFJQC750s9aGzl+eGPCKr9rsTkvmo05I4ns6Qjh9kOiVPb
vZseAbDpFjepYp/g9WHLyPsD8gWrL98JKNZ4QzcNohm9U3fYlBqlYGc66EKu9lhlidSEBmDhUS5W
kXUEcSUSHzee51DLkkODuENwlCvy5qm9J2Px/e7WiyDx+bdzZ5UA3Qo4BqSYIxG6i/DfyIF4okHX
eDHXDlW8vWngyIZBSYgKv3scJBDzbBTsfn2LnTtFMKwtw0WUuIqZah2fkrNQEF/aPb1RB7eDGOUe
sNEMhT3nNjof2q+pY6TsU4F2xReuwPQLq5vvElHeS/KnR1Cnd6NrZlN/XwCoqd67dBOdVcd3jzbL
UHH94KBJBYfOUxHi0w+VhGQPLrfzpRHoTyt33wrH5xMH1OaZLDy1+6NQE1ZlHOnPM7DVuO8zXbUR
UazfDvtuzQHr0fPpITYecPb7TBEIFhKquSm6ymD8/RqJQ1qZCSm5UgCkjttfDz9xBmShWvcvujC8
EbsrY1Vs8bze6kRU/Z5ryikmkcfh5XkefUPmQoXVRPWspobhoDx5bB3xdZw07RYpTHrSj5SbSnGt
ocFyqnqnvxMRVY5FrCyIaWtCP6V8e0qrWRINExckTqxGi+ChhB9Awjx3piMF8jMsVIjmRpd5Vmc9
3wlwzJVo9RdmhbODXbqSp00bvxON4AQ9Imc4NvoKja32z+xBV7A9TXNQjWJvaOIPeb2g0SvSaf1y
Hws7BNsiotIro/SvbCyGPieWoeGS7bAG33rBYLuq6IMwDGNbI6wxLvRJ4INhbyegfBDX/IuMvByD
J1wmPTGyjdK+JnxbuM0+7kkIx2IxJZPbDCTv0Ryznf2ZH2M4Nqbv3+JaEcAHPis6sewX6c6+h5/+
OV6kGW4marlu0ypzoJ/v+Zs4NnOlIEUbNN8TyJiYmcvO1ok9punUCzA8ppXII/DvLPMjujP938OM
tiDGOokx9S9ZxrC6m3QB+bVP8wOZz1qNcmGO24EzFM7FLMwI89TSs3zRStiSd+IJ4y/cBMdNK8cR
z8cnBVYC/nv5+Kf1+1BWBoq5crcVPnOHYvr8QYzXjq/H97peUJfF4KY5Q93riLDc8c6WkcEkIVve
WYiqVjp+tV2w1xZ97lZ8xEwOna1XOhtPeNplVQqiFcPi0y3r+BRziXkLeuAebVEclXsr1OGYK4Ym
961+OPZv7qL+wylhe/Po2SmzbkXeVZtz+En/e4h1lCUcpvmd0Pqo3/5spzozi3bW4cVnTh7NhVfC
+V3W8tbR+LtsI9IaaJCIJ0QFisSTdsoJpoDDl25kXkrfRzAEXtRVzbcoZr40onvrLJKPE3IaXYeC
oSWYxwUhlbEbI3tzUg3No5Hbp4juCCyuCXsJUnKtoWyR6mB323mrr+8JHtaTWCLYFBsD4RVjl4/2
BGaKYwXDiUQk4/ppWxBfKCbmuk2jZMOvVGfbGjTc/BHR8w+yTLIB7X2GLfjE9oXXHiaGJzwsHGXn
Qt84S7K1etM83O87pNZKCYtGKPFYPyjo+pXK6BxXFTnt51PxCeFBwFPD3X/anKJDBXRHQbcWC+4r
xIm+zPzsPky/MgkShJgor/FfCDIa+wqbfHJSeqPe5Snm8YLg4VS45c0j5BYqjhDXiw8lFb6gEgEK
DW3mleFAfoqtMRp4XH8JNpmUpTzm3aMmPucxDTZr0jXHDM25Mz6OEj0MqvvfAEdx0BTdIu/oeI0c
Y4Xf4VRkF47B1AX5NVUuDHE16s3SWZYD32szsUZh94UsWkuCi8NYoZFXpvQnmd5Fcrv24DTXb6uc
OAb/POo24M6xqdKACQuqv1eVdAIPjocj8zzvdtdSzGwtaN2LFEpEC2O9VfZ6hyZQGCdT0fz6j9QL
b2V2d8j+GDa7CV6nJzM4ztZzHDWVTfDk37rNy8y586UWjm9yhyvPU2vCqx6p7Gw/PUsLfooo9bYi
oKeTrEfn452SxY5of0rMqPF5TfbrRkmwOgyW1gXw3Mev1JhZZ3Ue1Vdy8Nso4dfYn0yFYhwoGJpZ
8JywQoiqj6rPR8+wsteNdPWB6Zt9vaOS9B20WJ1bU9xQ4+/WF3ZV8cVScPeHUsU1pZsa03IUpZ5q
T2SNnAWI0S3xkVkE25Md/Amzf9pcGFK4eYuk+XY9bfWPo3CcK76mjl7B7l1KOfTOqX+GKSrVE+Zt
kgP2wnHPSXjEAOAbj+x/pFF/L4CgiY3X71B4QTjnWAbmvq9xf1ZGxpx1ttXdJhE04dXbwuiaeh59
JDqTt7QUPC3oRPkX9gxvc02o1KnUdZrtSNp8dxkITy8r9U2pGug0M5WRc6NnAABY7qteQCl9YYFj
8W7mQ0aF+GBTbn4eKwdXD3EOFZojIxCR54oBI3cZn/JK+o0m/yVNMzE+o8ZhY6ZkNYZbLthcZOUY
lEOxZC6ZGQk/NRn74/pMwnAPazJzRMJAxI/a0KQWckF/CpcsUxLgiHMJKNhrkU+VXJZjxju8W9Gp
GUV2Kxt71ol4AvMGaHICV6UXAt0x7FbfKy+zFIZGPB+ra6VfqM5QhrJcdgb8dFIV4cxQpVjR9xW8
YFS+o3s32FJSR836d9aeCWMvrHv/y1pKo3dFy/wSyUR/Vvnz1xOOaS1eQ6HznsCAsXC2fg9I/hH7
g7Zgu1HECAXJF1D53H2BUApCUpReeKs29ZngSm4R2iWvrR6kQJgdr/1HAPk36ZDAtjErde5CwY6d
/4TLuDkiWDNKGOI4MPaflKGxKBkORRZxe2hh/7trbNd9lqVshk8TftQN1DmNNMSDrgMcB+Hr+a/K
bRgLLgfqHxLFPnklRoGZyJeABu6fM0n1VheM5RyO2qmJOPbq6mo3mwm2TnIwqgkCX+z1l7KMlu5a
YtgKdeVFrD0c0tR4D1fkj919WrVjLCAfu2Z5Tp1RrC/wohPbI31TTQHUwda5WwqnNt1isyRAkeCe
bmRF66igUBbXjiV4/1SikRy10X75Eek0hjZJ7HA+/XFDtO10hv1ymVB0HPTmBze6Ti6FopRZddsj
fBCXDKYklOkclZiqA3fa4UpHgw6IfUCGf96b5r6PpvqTougAJwtJEpLHMEZxLZOJOzj7TCwp13Ov
c2Up5kUHYDba8dReMizKAy3oCPXkPFNVZzDMOlYgf1wj9VMnBfLH93xFIBpoEfvud54O2MK7DD8E
kn86rLlK4xmDSAYu+Jf0E9Sb3RSEbl2uB0LWaZ8MdN/DPuO/yRePf9tfgmGtTSPnklZJ388R1FBb
UaB0O3pG+JeoELhLpx6/hhK7iWHyZyLwzFOlUOidRFwzmquZvKUruADuyHdsf/flTPGz9zWG2Pou
8TgHcKNiocfcfzpuagaXKr35poIvRJiDH8lOzOvI0fzCircPkGkkblcY4jxwvbx6ksrXjEbBJWB/
pgnhBO95kpjZL/gEK6s/csSAGpQOyRxsv7F7m2NlI7eAdCQMIl51x8m/zMxE6FxSmtjH5LhTSnOC
qD773GKT3/jFo6k2hqG6bNp1yvvHzzp9snylaot76Zk6ZZTN8eM8dWHYaGqYVIpD/jOigkYQ1wMn
Zxa8DxQ1L0ou1icsm9l+chUeimzJljs25wgUQSqgmd10kdTpBv9TSgb/QtW/03FO2CHEz0dnbtcz
CaKVgMKmbCsSz1btVXzzOsVJuJ14AJs6+rXZW2/b1vVteFoapDAyBAMrpbyMM1M4dkjtmbbWH2ZW
Tijep1vCnaWiKdhiOOW+ljSmIg+qzfGNxgDsjRTidfOixxIIHU29f3dWRwGg/HkNIzgk0uDSwzIa
xdqa00gstmGNTIzGCdg4tMYFdliD01k7xybHNugy9AIUUrbTc8vuSQrMqSh775tJnq8s2u8KF+IT
ITDzzdU1WmPBMxsBUF/wjYkOmY+NEG9cvZSdwAlhJRjW0P8RjlrrmwgonXDhXd1VzwBewvjiey+V
PyFJMqcLW8wCiFOfWg4OPwQ1FELR0F2USPnSkjvcen6vienDjg+ljP+y5YbW6+iNbquINI8nVbrj
Xo55YX2DMD3leWQEjirpbh8u9IQz0im8lE27Bvh31RYTctdlvDQcZDwrIvJUPHprqYdaZGeSDkJh
7aHyBmXGFo7yzqllYRAAd+WST+/LcKhq8v3x+diMYe1eeZu2dLp4c5R6nO5HkcfUuGKy7QgMzuDz
QAiEENUtf9dsmxJWUMM6P/m3U5mSzYotBxTPOXs/vtvdJBbkpBU60NkERUi3aSzGrt5Rq8bHoKN0
HzxfuUxb5W3R2NU7wb1n5mYh/rRJpzUKwBt3VVfcmBAUDDRncsYlCcUfFHmIXFrVizqnXmP0q8ta
heflVTqjTSjKxUyNxN+/luBZkaNx3JLrDWK5USMVAoktL8lRJzOXRDbZQiwGajbvrPzKg/2HMS8O
KM87FqesFxnBMwx+xmNskP7rn1R6nJVY0jDElgMkZdPwt7luruea+hA4OLfyxalFuKjxRqmPG5oD
QKsDG0TFgd1voxMhLBibUVGf3SAUvFK4v219Ek4Tx8kK6IaP4ryBsWfKWddLIgyXV2gKtJtJo3ZI
zviL2H1mg6Yg2B9FYwRPWfJkhXtVz3H+fN5/t5JUOklF4iRPhocxkegvU8Bvw6Nq40FIZJlwfIvf
WD/fOSlThlvf1NQNQ2UjGE+T8tX0iMZRy00bRaFAF/OEYvtrb+mMUDWAg8hbDG+EQAQV4hXfkTxd
neoPGsTWigKZfUJv79CAMe58JtqrIiKl+w6QeAmVFA2a2UhLv61kOESQKmooKjANCoOvvnE1Og4T
65Q9cTPosFLpajIvo3ytjfFCVvYMRcjITqr82UgH2xjB+UZqw7JAupuRha1yx7oAlJPPDXzqpgQq
0eFSbwnCgMr0oJqTapIm64WUx1KKDChCyN551twbGZvRaMMf/io6uOSJvbCuopc4YHrE9FPNlsQQ
X1QcDKV7+u6a2TN3YfphQjZGKeY1gLFpvp6p+r5MPvobhYiCurNM1qD97zqBaNh1r4oSx1+aEyWE
JP7d0Axo34WZQvs5yuxbxXXvUf4gegPS/85rOO665Er1Yvo/z2TfLbvmeDAMH1xbsvQRyx+WVys3
6OuB09FOZmMAVcHDD4VjGURc0cOKMn9vmIDJbLpXQywfaN5B+XVk1CNSNRM476bgyIBd9Yqxxte+
TdPiTsYjQxu7MrpZ7ptN/iZNhiEEoF1Uto6S3TcnY17pwMqgdVxdvqfCeUyrJw/plcWMnopY9xaL
7JMeF4eeYqOeJ4Xr7Uxen5k87y3szx0wpPedtIOUqj9U1Aa6FBJnspwZRSKlq9h4mxJzC6DsLo2r
pEvwVFW2PS+jt/cHw6Vr9Y4PLlyHiyoVD0/cV3Ut4WdeORG8LZzOIHxezU0z/LJGDMa/27aERaA4
vBd2PlT/1KgjTOuXwRh0qbirzaEAfRvTmJxyzMiYoi2d0B7bsRe4jWxJfDvJEVhN56MhXZ3QlYi9
eGatygHB8hyKmuRJ81BW47Aj20tMQ58R/se2F1fXzCBPAF/rHHhoDZNVxojGyncfERq1pfcQ7Tj/
K4j/3sUKPECtFW/gKsDhixXRxSv/u1T3AX/rxbZBW7JcSa1csjo8L3dkiDd3orelHQ4DGAPZfyHp
9ca3ToUP0xLyHqnwJwvG2/LYmqWUwHY/79BFoylJ5HO63BcpuJui7gr09QJySiH/i5q+ntxWZ7OD
/f+YYWqwlXasjyATAI/Og03Mf6eHpAO/A4DYiega2zlV0eOKzCDWfKRMPGjxh75/+J+M3Z+L2w1k
0zfSAT5U2mCfxA3AdfJpEbUPqwUxvNzpOBFzWSOM9GVgZTTJYx+FlZAserV3ypQchvonh1HFI7uC
oMgipLsyAehAEhCYlaP36B/juWo57JMkEhRGj5wu5gPs1wfZc+5NRGOoLCS8hynQytOz6d8Y+ubc
DPTZjbLcP3x7hKhq+1oX/oYuHxiCEBqB5J9D94MPk9VBdcLWoWOvNOrIx2DoiM7aPRkOtsEtWqyw
jY1sQ7ibWBOsBCxoyPtLb1vwGzLuZ3jS8SlZQQrpuPd1Z5chu+Xxeynweytg/H5WA8iq1kyus322
J8nhMnTZzbrNBC4oLBNeUruCDn/P3mQ/YH8PxNp5N4pbjpJbe24QI/akBckyNB9MIXpqf/pz98tr
w8TtcEAF09cKA1pYF+9xRW7hygLrtk+yGPaBgldYBV9xOdz5fodsTVb6ikJPSUJPq+YjKewHd2Z5
g26CqWienycEiUlVpqYAnkQXc1uu1fzdUDHqmd61L7rFMd+hBLq+fP+Nwv3AcT/3irDXUNYTcwsc
QFbNJgVJH1lJxCkD6ZZgHBVbMt6RCTSkVsC7QZxFQ16G70Cx+LxqhG14Rtsi1s26ggc/CD4tknCI
qcwigTFf+iiFPF0oGB7iQn/wOoG8MFRhhzDyr+qmcJ0e9qb1KMqHNqKv++W4wipX1Ivb4OpL7l/W
03DoT9FX7zgZzZd/zdOpQaKOnb2cOFKkY1fN3ysN+AEIfnOTxSL0jS+zof1tB0XhEduHvFOFn9+3
UVXKtd7WmF+BYzS27j0hDQ5YjCwZpH7BJ3WdzVT2f8AiVSdzX40Ctt2PC6OqE6GesA7wPXReD5qG
LqMgghb6jusHoAheBw+UfRJID+jG0T7/JQrf6xJjUblWbDK5UHmnG3XqSgA2lT3sTSTCpjwMVJX0
EZhQeLy4iahNDDRKlWZQK5iu5D0jbcRThp5LPVZ8tHLnzTEVpEUPzXahSMuL59hbA3e+zqkbxVsI
1Z3jaQCNUQslpiu60YkZIte2ev0TQRZK184dDKVW0v3QYLNEN/GlYWEPTMDbBSn2hx/7f6VLFQc7
cyhU4Lw+6WVE7edD8EAGQ0UYuOeMj9Shbtv4Ed9Her9+yOP6ynFDUx/7au51JKr9ACcbHkgrBHuE
ND5IEIJJjJMKp3viEw1PyD6/jNb8fK6UziXiqWW40pD8C/ZIWlA54c1WqmLQdc8UxY5+NR/ptZpB
itMIpHSY5k+nQd/WspW0AuojxrsfJZk1OGjsvSZFxX0cTEwappcP4fPcDIscYX07JbUog+de+/l0
bpOH+WOPrNINNKWTvcqeMPLeRoztfgIIxf9Fx1W2p+AZfB4QweRdJOZ+yHRiHFgWBWnsXMi0LLZx
WHhnr5qj68jZIQZkniGYf/+WeG1udWhfWH5Z83VyBoUcHZi628doqJg4RcrYsnK4c7G3GItt8sh5
/r/u3JOd7QcK3W84EGbcn3/Dr7CbQG9vmAuQwUczo4XEYd1nkxQBq7Lo+mhHRnvSyqOoQu0uiN2P
cKA6yn3njsihK/nlG/BF4PHNtqLUgWOl+5ppiw4LPBR6XU9UV/SCFQ2LHw80vZJbVtEUcsNMxCFZ
yglEsXJ+A11VPF1P/La/Vk0F9jejOfTMHG9bobJyj2K/L9l+Me966k//P12UvtiQwur+2CI04EMf
EJ234c9+wCGvOGd0pUi91XAHMAVV65UY63GVvWf/3Fc96J4NpjI0t3Lh+heTy5O956B/ee+jlDIi
uYfoTGNEEqG0EloxStyv3J5rH497MIFy5Z/3GQswhaL04fmsDt3oSv7MYeTwzD0aCVxRNmcED6AK
JNEdyHegWMnQM4TSERu/UvwenNtJGCUHoj1JDXDLNkQOs/DGzcUFZXlYtTBINzyI6MqZVqNcjMdZ
vLdoBMfOX8xEwf/fR9OHyk3ZEYSkKUw8Bu8yUXPFHT6cuOYmkElrE4K6d3Mh45t6wlFfnjYX/p5B
tUYVA7fSBB+vxCJlTqzyAbOjNFXBJzQs4P/jlw2vyhW8Bo2/BtLWzzun6X5ms8d6Rbtwx0CHKXNJ
E3qO2xB7kk7Rwpro98z+/8MgaGOV1K5RB2bf7hcd/Q8VIKslTuSax6FnMDDun7AndJwOw49EqPwe
aW4Tlu+JTvfDe/IovKhGZ+UMt9INvrRX298ZX85geSMlciWGQ9F93aTUnOZzF4G5gcWrG63ISo6Y
uwFmzZYTLZYWxWl40fpKOTTR7EZc22XHF/jCV8i6Yfq221dF6crzsvBx50he/ltfTloYThohIK+Q
LtCH58FfiZEm+XYm3Ew9TGQCeBglbc/KjyouA3VReXzMeVn/g2JLEINAg3POpRHMKp2eUB0lUW29
dYLm07KtcggIFeDxkWn9vUTdEqze1IWGanO/XJCVYFkrLvOwG5xd+afZG96miHp1K38QAFUJ+ldA
2i7dOQm18jWgvLUY4Xn2cfuUUVgQ6pqz/kiK0u4tT6kIrlFZgmxDaz2idpFR2ZdBZCfR10oMX1nI
3+uEWPDmauA19tFUQzEcmTnkT4kyz4H7EVnyLV7IMeYB62EsH1noYQA5LQED/mRJLVEeo/KQlbLo
aghaMMXgVJeWgtmp/njFgxHT5hqYhhWRvWl6cxCHS6ttaMyhRRgoe3wYIwcw60eMQALd8w7G1P7F
4+0uzPRsrZjOimupu0ZPvm8GPzNxnnrXsL5HpADRtGQfl8mMEKoLT4zuB0UwFm3V6b5ms+BNvEe6
pYVlmDEQojIoIZ9h3KL04uUM6BlDd95c4o6l377+B90cj6PpZR8MepBM8XeigsQhM4X1HvLm1De3
V0FrSj+ErRsrSFF7oM7Z1YR3CLx9guPHO1mBzdukpipmU3F9C7u/XGM19wvYkp56qsQG4QGyOp5Q
In0OUQqvjSKtH3LTR+2gVtpxNAd8QbJ57QucYp/PXyvsPM3uIm1VcbzAq7vHkfHuRa/lW3pYIW3+
MVsglaVn/+gMZT4DS0o50NHnOPZmmNrEtdd259gm3F1l9j/JfRWs7A66W9DFN+AGwefTwQt3zpIV
Ml11Y9k1+WZ/2nHsd7NB/XdmGFEENmdcUOTV9lrD88t58tBgCFUwdFancRMBURrKxtKyGUvBzJKa
dhKv0HR5tZf+o/oznzup/baWYbTYqikpozGSGEbfPj3hHlcaITlQOfB/ZizVFneGBLn3BVPKQTQt
Y6DzpPYlCCbwkycYyZVzXGqUalu0W5nOE9lI4dhgiEAKzeGtzBILi7y6a5DmS1DhavjTajNsNJHL
Hkw++Cwu3VXELG7NiDL0r23dkXrzPAPI8+awBwUSrntfDw4zfqay/xi+ua9E0LENFqjKumCaFO5C
KJSeXu7+OkD6xqg8tyxLy0nZUbwzHSk0UWdAJ+dGz2bFRhah8Xvfz4T19RS6HEbTVuKOXft29OgU
CgFGd0hKXqKQtSg0HsjV9NE3Io0pM73pjCuJeJAPX47AxUt9idpMCxz7ATSj8QMM58c1OhVjFWNy
iBehG/uxqbuFlEDPEw6TYT6rPJ6uMMYPNPDs6nkuloSdTNuHs+YILnj6HrZEMelXezAzR3VHJvI+
l920QzIoa5FIXBQLT+i5NH2gRtRJpKGRF3Rq9/D8oRK08nL/vYiHgeFUwCDKzVvX13HYRm6Ew+NY
/CrFOOSR4m09NvgY8/FX1YV41uvghCGhQyt9vWe5gDM49nlqqi+pPr/WVUoMcpp5GJv4uiAL3IkH
wPRIkNrs5wvXUnPmD1GK62fhvgu2cpaRkEm+codAQpyyzR5HStqqtD+x5vYuIj00j6X9FDKv9GBa
gc/5jlxbTFwHIyh0CggCkNjrU3w1LMn9ChGT2UoloSkGqF4ji1wiAqn2YT6zSLOfYXKhFsKUKxsG
M7l38h23rAM160ssAT9kPnvIeYXnsTSJijO0pm+AYDiSsQ9qImoX0f7PWb5nTzlsb/EhT46Ep/FQ
aLOrXdm/WiBejywhZ8LTnaONjXtZHF56Beto14Rd1WKj5RSBp9XjKmxR8DMgui1b5qYI5mcis5wB
VHaDyQbQ4WwVH21kXb4Q/3sf7yA7x2kEvF4tisJH5NzXTV6UCl8EsX8h3arBc2CE5vRvloX/hrwG
A3YLMOeqeCTM8P/sUIeTLvH2tuyd3lmf9LaL0aVlqKBhnTHquCI6GuseuzkUQOYB1VlXbdIR1C91
gVFXUXwcotlyFWUKEZIruCiiPJ/x8xMtC0YcpidzcNgZNU83LWBgexJsg+pdIxn0DipiUXuRBbe+
8PFfzj5SgZo5bzzw1ig5bw6DNnzQoTzZaV2nfUA22/Lzy6E9Iljye0Jutlvo2Np5QFrKkK6uXRsA
JqkWpqkZD0yC3zL6Ufi8wsmpRy9/wW3jEnFdHeZ9lUX8AEBnxtFxwF6j3Tl8nJNPiyW1uj3z3Ga/
tY8PUG7iT37xJG04Trc0504ZYFajkf4MXkDcDDT2fkhEF46vCoW4cRHWPpshzuu1i/MbggyjLI7g
zJnwmfHXcWX1TlFQZhbC0ZxLUa7rXRk8ICkQz+PnJI8cKjE/E2A24LjCvGGN2so1cQRAV8AbN052
EQ5RItapddX0kxaB+3ehJ3mFRYsDqloi0WliV0FNCUvvzy6pdLbb033JXLUELpjbOVI6LpE6RqCq
eq/tJwTGy0I9A9wDcUtva6jSmkqpi8mAVw/utLEZpZXjqTAFCmk5sddwxYdGiBIOHwFZFM5hS5kM
2HjKokLcpmULJEMZmXPM4zfVenppOy/ycmHQ3eaRbcDOxQg1C4w1RFtuuHnA9hBKYuUngTT5LRW0
xDIt60a36lZCUgi1Q5pX5tQRpI4I4fkIarXJ38gd8kbSRUfrpRQ1RdqTztIo2hOiYzGaCtUtZjDz
jpzsmZUjbbRT5e43SVND+DQjMz/Um2vxjBWvGzRxXRKNSR8gnOTyHvEG6XLhF+mlwzgXBECjfxJl
MxVee+5hES4nMyhiplt4r1/tIKUxaun12/KOAxNdIrNWG6jfewRxO0OdLIlrANrYiaKJJ+P2pHoX
bI9sIafzJpjlI1opNq8HhBIe8QxDEvmbWHx4/5F0Vj03NYLEn9a43pOKeYivXYnuACd4fIAohRPX
KSGuIgwBXYhSVgvn0lsTXFLSb847+mmjQcMsUGyEK5QSYWMxr2sVKh8SqiZSCcaLL5UQKaoL/BdM
u7lgOkuiGSIII5XEzh2Nh83TTfXgtNlcE/FRBxS03S6Rp2KqM6GNTiUKcdsdjzwmfRKaEO4gCB3v
BQIoLr7qRGeZ9deWt5Go0gbVrUJ0dKDBGNMeLu+nbbA3qK+Re2CS8VwSLSh7Q5PmTckKjBKcCxmc
ujFHoPkvGfP5d5xAaynRE3oDyLQ/4S7t2pDBl21CBRtKRW9cHgDACFhDnFQ1BL0mETBwvT6oXE8K
qntcnqWpTG9CLc636PqrtT7i7Fg+8/3J8WF1Lc/8jERwIV2c3S1xjIHzFSr8zyJ0zOrrCUMPIMYM
kty0pE7m7z4n/9IXgXYQTqMVjpZ9ODO5/mjy7eium3xL9ci6tBpXdAb907tA85REKg9o0r2zAITw
a8qou3wwf5qlvBeXYR/1VEzcAB6xk4SLE0e6ZCXsVrnMD4RnD0Q5t6MnQ9rjIZfCCExkSrBbS1fq
DRTWZW1oGU1KrbqtzWRlpA9k0IinjJcEM+hZWfuWe3iSPE59B4fiLvO0iZ2vVIYyGqWf0xRQ6Tto
0gpZH4Nr5V07/H1L6ptIbFDCFqDnBs2m3JzvwxDcUI4MDiO2PPSJR3SZ+dm5rIYxfG+80oJyqVS/
2qiZQCKiU8r54LmnpmjbXtg3jv+EUU5c/pK01mhgKlChRjNX6ScbRWdxL8ZV8LRTBCp5pTOse5zY
daJOWvH/GtgL5p8BX2LPti0qtLokdTP9+7AS5PLa1oLj+Jag4ivYCGyvc6nmJUS4lk2N44em6Km5
7u6N/CIeQRHmsXss7syL5iUkq7w6Aq1B3TEtDkApSGTZtborDWRi73sH6lrSHfdJNt1Wvn8/gh4e
tNiAOpKlc5tfC+G7lYXkiz+RerGfTzj8BGzGDD0+XIwuWdV/8ds7Oy+V6LbIyykK62YzM6yM/v2/
rdaA2CSJThaHWdUj8tTA4IRX5wwBebLRQUwqtAKEcIrXRuVVmuyXWns+r+D7ZclYBBnF2otrfVdP
sj3vp5CjBYPYgGFvonC/Kk63KjvPOYgvtMmORZ0gUo71d71+8kcaTGScxb6hXmw36Dz6tOXHVOYY
/IjcpvyIg8bGTOH8tquM3cjumxPdQqE0vSpQxBlns93ozAvWk18x7GnRomHUDGx7AleFzZkHjyVC
BmlCXggcgsg3YG9wc+Aq40S3PCh7isCwNWj2er/pZr+Dp/bys0TzA0f/ZCs5ExY8AJq64ySOE/Fy
qbsfusl5+YojSlyzuodMhYzw81bAA0eB0I5DrqOLlCYEuevIMGOGP7JcIHrVVi4NLcXV+ic343+7
of6FV4sF/07oeuULMRKNncYCkPgrsstohITWKHPxixnoRIDtP08hCzMGAR5Baq9QwjZd61C/ARXF
Bk2un8AxOWkMT1gQ20aZgx3sJ7hTz+t5ym5dwwW+oIdSKPOVjSzJcfGCEnEyCBrnIadjUIgJ/AK7
kZ663rS0rBf5natgvSiVXg14Qf3Pasyb6X+fZ0lQssm14kLfUeph3Raz2qymG/NsdxhwaXMGlnQv
oUxQKNCHPBWvhH9TiqtKr08LB/K0QX2Q0cH1fl5PYRf706yisfW7ui+SXBHb+6VQHLA06lLbHRzl
xRXyozVjz1HaNR6qrRJsIAb2WtjZkq+0tZyvaHW9+335KVmHfoTyvb1UOIls/xfXsz5rZcJ2wT7n
SiMt7VNCDfCcaWsSAjps24QS6BI6oyp68qX5vb6kxx2fZZ3zyMhuculx53jh8fDLaqxBu4Pu9s+U
uuBxmmmYXHemyuW5QXgrd7jZLzzAD8+0Yzf8+IDLz/lD2U9hfNP6T0OJMIu2zzw9hmf+V1Ael8rC
clxiFWgegmP9o1nKOv8WKss3gFq2NLmYNuSYMQNbqFZw+Br7n2fDMTirlm86cH3HS1qNM18cNNij
7ff1iTiiVVI8UdHEN9U4MHZEW6dkD9hX/lNc1nK6f8EwfTXWzkDT5azX0XcmjjUWL1NXHCqlHDi7
lnjgkrq5dztJPF6oBYwCdbA4UT0nbMmdBKkB/1RdylRjlquTGWDNIXXXzhnGyJaoTr6RDMTrGH7B
Pm90DGOSQ2cztuwcXHTgzMwhLxoD9nV20hKoi9imGU7tw04y5G1lXxPhkMYsDbFrEKojnBJbWYBz
fRI0BXmO3yFEpaHINOzU11pPGXqtl/zT/XelsKx33ofTa6Z4sNGVyrFzRbceHjI+XEAKms3anzCd
p019cHMeioSCl6wGQdRuCM5k3PdAhWhCrhm8k/ABczYOHypofz+ocnUhlRPUNh2oUoucnB2/vaza
Okdq8B7ibBXe7hbjoQDT6UdlVDh5agYBbwMkxCNTDJnu6P54PhxVCrRMU+B8YW53KeHMG56pLEOZ
864yUsssR0guY4S1Aj99yRMb5TWxmLjV97xbcc9WbU4Au4T2+Y8KWgGW+NhaMRElhukReD94+oAp
qyi5mtKm+CyOZ0WNVaB4l9CotoMu/tRiQPX68W+X/ByNGY4AnqXJ/DqJFrPjtbXySgoegJViHEXE
DTDr4UWq7FkhwgbUj3MbYdqQDgzg2IQ4GllBYBzsnFHoeQRI+rNrWsCPQa3C/quFvQAqmY1WfYUP
wN3Kcmu7Omr6J1h1YUufw/t6qFlBlCHOTv90SqcJXgNIaJMooZ1Dt6DHKpvBASQpTUo7r3gRGBX5
3OQf9hH2Rr9q3/egPXBUqFPMqRnHJ4M+UF561n1MX3rM8O8EmUs4d1WJmhvHFRWWH/Se3yV1Jq/z
q0+Rc2BsBClZAHxbQW7B5Be5gggyif04jUdiKrnJfQY1fQB5N/W6ykQ828J2IL72t1Q57IIa8p4K
HjpFChaBPcD2MIbfFrW8dy8QlKsn+mXp6X8XeFyWrscGzZ4SVatA+aeBC8qC5I/WEr1+Xa3XtlpA
HSF/g+IRJQ90HRzBx47toS08/Ks0JSrKyrP4I6P3rz5geFsRlavViX2dmQmvxmW5llmoaK7mINSi
sxzWOhHhzhepK5wKLeyg1jqM1ekhpxW+OgF4N/42X87nn6gdN54ugjLL/pbOzmxtSyB6KynoGsLl
7/Kn7dxVCXIFNEGCwPAn28VAuTxelE4xSuT/lZdMjoXlao/CKxjGL/2kNstY9iZiZUKpevciSGGL
n9igOHWMhKp5QoBeLaPwzSbqV7rpDF7s0bQDocUCtsCNOsvw5Ms4lWkrprLdqLCjmAZFfPpjjEA8
bsfF/kT4+QQLhtNHtoEpJLak4hO5M6vfHzXMZk3VgrAEo/n9RWSliAZOn8IfU72i3+w+I5TSCaYe
gEknItRsL8r3/AEqwz//ysLJ0QZM2y9k6RjctjdJ86WcA+D8N/ViHPBCjS8jpxCT48dUDyqaH1yE
FjxB+Np/rd91SqKL8QTFnZjAZLJu2PGpCSICOno6m0UOktG076KexFi9+x/UOZ/leUslkhXlBCgQ
W3RIMv/UyjB4tPdcQsKV+VbxrsUQYyX0aU3YWgkyIT6UscPFhPBAcqNMeI//IogZw75gTNVXrNAt
+gm2kHQ6Iqc2taZFwzUkPmYpnGlfzsSzGWCLm8cuovdH0LI6KhuvBBU6yUiq/oU+zto9yRabFTFa
B3/XldvBwnQMDjRt2msyhE9OYn5ASGFESt+mXXgQkFlCv4hPTk0+spxkTct8nldUQnk5zMgRr/+k
FY09bVI3u5qcMS2OpiRVWqGTQ3xQcIvwAHrBTTqSX4Bui7Iz34HDzKcGCInISDLAnRj0OHFo1shX
i6WKQSWe2B/5umtS1PmmT18rKbE+CITbBhBYKQQJ+w+0zlOmXOoh9sraEAtBffGg8fP4ESkHbEcq
vMdPQ/ndMImfmz+pDAqcgCUJyAuCH9gX43kE7Bf4JwwfWeWeHNwh6pt67OEh2xE+qke1AHTAnM7I
M/3ig2nbvsij/1LFruh7BEGm4pl4kfco54WNRjECocf26A/vrdKwdqWRYr7hl3nVw2eligUkqb5V
uDBnszPeZcYU42Qf9bX+I0PolGAN/HigvElyd8jaLmVHtcPy4yqcwGyP5RaymyjfS4Pk1UOYtjNk
fEtiXPCqgzKzFIAPutXBvhVAJ1g6Us0qtVfgataTc4QqzDBsKI3HNj4b6vjqOXbR7P7JrtZzZ39u
0sKDczs08tk8IYFjqLkKKkpEB+TR+GJZdO4pcrEkeOSMishUlAJbYRu9WflaWAaXBC+V9qnPeM3e
SJNRKmXQZ6y1UKHYekVeJjUpZpBym2gaal0m0B2HE/FgAsdyvbfLhsNKHGEmyfO72sd5yzopcc2m
XTx6PSDmXUVdOGWRRNaT/K62hUROilnrHKwy8gITvcpj3mwESxR3w4jR9byVQPs7y2FQvRNtyCwK
m6BQuLhlTQ69ZlY6AmfOFxxOzmLfWjs3Uw5cFT7drWiV+pJyRqqzRlny6xxnsQyiwr+sXsRncGBF
/aXhc17GKXkU3YBkJ8uCYPsQyLpFQdAIvtb8frAp7huh00YARBr+QkhMdHiLXIKJOphZviDjhWIs
mZ3OzaOlqijBTaQfsNA4UHCtX2vjPknMzipYyzC5SHqVdtHDs0IMTAfmlr9/wAMrs6UhqL77QbOk
zYYr2lPSQh6BxB7mYps4b2ivR8nZQZPmXqhj6FErUGKEAveIhtUCLAqIgKe9zcxqyTBzTQnwlAeS
N5VWOnNXB9MFS5F3AFO2W/TJhyGAdSf2zrDalOcykgl/luSNGzgYTbw/VQCuM2inu2jtwUwppvvP
sN/a7Tky+yocvAMr2h/B76PqdTZuCD9zcSWaeIVLYc+lzQtd6vSy6yxBOSZ/fhMPNV/AK0y8s0fL
3auVschqJFcIgQy/eFoN/4l7L4ui/jcl57hej1YDV0fglln0HqmQv/ubHdt1GT2vnxreOFiQZ7zr
xR13SJntKaUxM1OaDdybj/m2ZRC9fvAGwhNdql0+4uRJGQ2nuffY1wqIe+8PM5u41m9Fq6aZjbKF
YVIpqt4M3z/ljPDkhdKK+5RaXV/CTPDrE4w29kw79U2KZE3BniidG7Lc+48sfncjTM8hZ4ujkEDm
KjNLKJpySI9EIPmbD8SABV9Cs0aF+tT4x6UQQV6YKlTyIwhRmlIryvjSfyKYUyHbwgEkEHAMQ4N8
IxI9zJWszYVsT9EglE9cOHtne3LKUDzW6Ahpa5nAzHLc3eszgHNQTlYF4u7g/r5aftGtqjRy8eop
Q1Xm+91kNvCehWNMofyDcFdzw0sPRQ9JMjGZkLoh1zicK3DzITYaewEz/ushz9nrkWPsH9UqWIYx
F1aAW/qMLh9GO620t2jDGBEBv+SVbBPNMgUFlBu4bKhWBrCzHFpmAWoBw3U49uPAjheIIxhQpbUL
SAH3cPnDVNhAYEJwyjdT/3OLpfsWDZ0CHBb/Gi2uEwhIVzRr3rYvs9M0tuQkVPPgYzqvuX5Of4xs
QbxTK08nvaX7lOctuBTWQ0pjYC+xaz+Hqf72QDspD0jb7BiuIY37n/qjzwc7GAkz1WPvW5qI/+m5
ZUPcOrDC6G6ygoWOa6MVHXnrMnEvBcnJWyVG8H+2g39PK3Ww0eS+sC0mugTlTwsnzbW1DhEtHcaT
1IECFCpXzDclzK3Kwh2Cg5MZJCf08wfRFs4JgrHIxSlcjWkar+3BGIN+lEz5rH5EYokQ2fYQjaxA
LTmmULzyQshKwuF0+g7t9eQVSMYH4aWR8uvN9jpZRMuUVwcONunhvCL+UJZFmub9G2dLOxe/OsM4
kwZj5VhJ/7A0SdUZVEwyvZyMqmWJZzwBDhJNeyMzDc+dYfqe15m5E34MRXMRZFFr7P5103tkXT3y
A4sR9WEz1kYiP1XxHJB+XOlmoScx80hqxix8meDC9aeXk1/t6EE4GL8gDOo8xwcVVRXmP+F8LPsX
3knJBwZDSkbEm4c1cd4CdvtWrq6lCTRfCHtXstjto7m8bT1OKPsVIAMKQQkyZFbWgoPsIxQeL5NE
HGTrrW3I+IfdTD9xNZlGsORSRo+nu8rLxSnNCRY7XkMUtc1uCwSGHsawwjgnhd9TC6JYGr8SdrdF
ATY9wp0beSJXPEAav5Q0yDa+LgCekeiKdH1AfWUBlzZaitomIbmqEhy47f+t2Y2lPx68NLScdENW
qeuGONPIc+BKyXlLMLj7p+7biKsPxkXpv73uNK2uRW9S5LB8hoYH36PncphrIMcMvNivutO7T5fl
8GFKZsGSsh3TKW5WpGwowA3jW6uvZOJsoYSACJuMvsqjCNyraWw/ZMwfTwAtK6pBQxUr4zt+IYRr
X86WjTivlUdeUdLK0micIs2eYZGcraLQlpg9X3i584z7ieRug9ndwdlzO9nfaSQnI2VwZ4JSbkIV
mqjaqs0F4OHc1N2VghIeYZxmB+hbsjuOOrItVqgf7XtnIrXb+s7g237K8JXvbHxY8rX+Yu7Ksjfq
y4TRJ7gdwrx5Q7jtYxR+IwvWYopS28CEDM0yTctZmP+U9+oSDqNaTt+mS4Se1cpqY12JBVNUO1TE
ZgxVdV/+P7m3ZtILiOU4+LQJEcTJbqeozUqLGDn/ayF6In7mbLvdjaZKtUqDJLIT65G/JlVgqJ8l
mTzbLNg8v9MkynmOe28jzVDdNi3fC3nbCFSGtYurPV+XxNeNdaVvBsDWvuf9CanYhS1YBB5cMHUw
47AYaHJjkjzbiWggufBctRrFjQY3WRdOXbRB3bcLzh1obl7EZ/aGcV1tzKkQwFc4T+HIQTF9G7An
cpiKUUxUwbt0igdLcdGzGcMJxDhA/ayCbichhQna/N0cNUNX3EprLqvuwSAVdOp8l1amz18z4UeP
Y7GqA6KjTabOSKq1Aqbquxyb8MHSghN9cfeuwO8ls3Nu88S216gJqfXZa7f8PSa2P5sB+3SlU0F9
kldIat3vr5lhEbO7xeESp96mW3avp2pn8g7U+NSB6D9LUubgbMWHy9yD7WAEFLwlqYfiyr67s+Z9
ZoG7FhIc4gcTgcFg9+z7rSKZF2H9MNA9ozqyRGntyPpD4eSYKciCqGAxKwSmuPCt/eTMjr5U+gUG
x9Cmxa49fTe2H6z0OX9+VtfajU/poZEngqLT3R56Wn8jhD3TSFx9eWBUI3kX8Xs/Og4WONWvtUkI
M9buxXSFJvQ2t2K3xOU41bv3+dNRfx5grwZuS27E5SkwzodeRK7VcRFW7rZPtM1OtPvbPnQT1zdW
rmSU6RP6Q3oWL+dyYdT2uUoK50KCX+Q55oIhW3B+EdtQJzJhOmF7xnJcAw+qg9I9LwerjXcCqSxZ
Y1snqadT++UzoMq5dICQD6CpfzTDJ0ulvc3t61XbeobOGy611MsyoQo2yo1+lGu7IE52qn5M343K
GOK+sW7DgL+7FEQ6hCfzeF45fFJx4wFfzFoKDCngJd3xZFBOP/Kd0jyI/uGb1J3eMpJZmcG3AETR
RuMuzfhC7X+SS9adIRn1qdEpW+lBs/H9M/B5I/kEaokdJVNPy5TjiD93m3WMeXTOZ6gn0FKXHqqC
GXY7ZAvGrGAGDwfy+zwFWqjcXA1bOs+07MPnvjPU/Vr3yCD7ftL4qYRqTIcMLWK4AfMYZSgJiHNm
vRP1lM5Q3EAa+2ME3bJNQoyAiFrSbef3isQ/fVJFTW7axXIemLwwTKdaSmOjd96/DSf/APfd3gKE
NKP3tPC5j2immxjfh2+n81W2Rtslifzr4xFtHcra4fuXx+lWBXZyXArIG4LAZyDFt3uMb8EFuUg/
+fhmo3TGKhkzTOgfPqoV/mRjI6vdODlU2rdlQtaRR26ry4okz+uyzHSga/OHdnvGC1IkkEf+iE5G
VbeEJHWS4VB4z1t2ef5xc01QMUrB2c31ADt2za1UGPAMlX/RE2mE3LbDdg4e7WPDgIcl+gmJH7Ft
k8ZkFXul7IvSLZDqAzjqcwcZzUyyQ4z198a1b6kp4HLXBYWRep0Pe5NqmEajbOeRjkyeAVlGx3bL
7b4KB2W9WDHDbVpedGnHQLml7FBxzZllcHD+gSdGtGwREskKhVtouZEYuZJsmnadJzNUHHu0ZD7w
ny0PhLsYa1ZeLBo8OAP5Mp3OWrs30pWaY4y8QPi53ZODlxgycmgg2ATi3zkGZGzcr0o/6icRGF39
43kpWi2gmVc91coOFcCkujfSX5L8IeqBlY8x8r8alMic6a6RHxKtc9l5B57WyifDaOp/KX94BCVD
/2zp9iLFe2MjhCZEYQ2IqUawYv/N0/QwF6TA8uxDLRe0LBMwGTx47C8mwBkN0tUjbVdMiHv8Cwbw
CWXhwU2qrC6wEy4N+wc2X6uMLXaJL47iETc4z4h9A12/nOAkmNfyzsJTLC8W3bPtw/YB7xSU3mx2
XpaurkarFJyrwnlOBptLj7Oslz4R0pzRuqLRAcBjRvgu2/FUKgxdt4jpH4MiiS3MuEQ5furWc55g
20QcBCARnaqWq/GqxDg3yG3THONHBVUJxq3j9FbpArK3llZHzNKo/9awf7Zcp2QkcwQAswLPMo8W
VtWCvjFpniYJ7+rk1kwpRWLiVsaygESj37i/ID8b4uiZsscgGe5nZRZIA0CZylv+6IlvuF6OywzT
Tj0yMcFo23ioeMrrMslXA+6rFh7pNXoZBWWqpBxKBcUK0a7TkyFi8gLkTbO3pWWurzsGsFqT7EIj
1bEfCjc42Xix/EO9xYdwLKexj0A8lNVjkV8FV66stEh6yAfsQG6AMv8ftF98pFi+nTXe9Yqru29p
hNzquoT8MyIh17tNrHdIwBrnWUk4j1IvrAf2v0iZYcmjCS5wHtzhb1XzX1JCpn5knwCxuFIxTEJ4
1l96BdhHix/CuC9UWyVDlYiFc5uqZGBAm8lR2nWD3RKutAGp2b5Mwj/5NCjZX3tG+uCEozIYztT1
jNM0nUQrvoJ6ilySDnHTcTBW/6s6k9eWq2jaIfCMM5gexk7Aa8qZ47/85f25bdUYboAzM74nEpx7
dxAUa+7SF/FZetd/BSqLxBVneDYK+dzJZ3yPfvjdmRH51p0ewSDgycsMs4YnDu+JKXUUgRyLnVzs
lSGfr1gGM8hOErqSzaxjFuuRbibqfFSo3ojFUjTcnNK5hNM+6EXRiRZORVRuKFv9mxaKNjw5yAie
wtfYAlGPskOr3IzB4uqFPjkHihycSYz8PO3ly858BeQKg+SLQ9+ZFJDm95POOziBFABMnUR3yZ5+
8WSWsKvwuZ7XFhHSzLFp64y3LMAGRy6bzV1iXs5Sm2kjzm9UTqp4bv3VOZ37+qjm1nZbIvuz3fyP
3IhJRmGq5VF1znluElmACy6sOWJBp6JAGuHRc90jpusuLb4T95SjspvL9N3OxCDaRFTkyCNcmsRA
nYrvCJJUuaw7GPNXkNnTJv82Dp2g5g6szTLDDz3y/FqalQCFgtsi8u/NBtu49hAqMZHRidgApv3/
K8L4MJSyMdifyqjxS3dLEC0Tig+GZBaErCPC65tuXJlHFIR+/NS/Stx4iRy5ncDNjTP9Oh90OyQT
qHfgAGizrNSsIFh5qFKIWB82tv4V/frgXyo5HjHq9Uzvdsh4UNXmjv7IjQCwjPxo2pA83AdR4ybj
/4aEddkjZyIDfYoBRWFYjzEGwV3udd4fDca0W254/f8pQ2FjPJn4gXZ7d4WoZswt19kR7jpXUMHi
98+mTFEevn2Y+infVymfiPALaa7AuOP1i2VPBfTnW7sD9UOgaMiD25xRBGf5FSWVukTmYTgFth/t
RGv09ORiB3t/1YDHMzg4IbKTNW4YTGOKSgVhKiNjBDEHdlasHE9KOVDlRjobi8Pj2BsxXldDORDh
Ohauosx/1D3DiIrARkuSFp0UGaYZFe3cc+nJFA6x5uraE1f72bCJp6gb0PilRCNPd3q471d8055+
b1rtG3/Q1E4lxlcu6wNbktX8n2BfFyvlQYHby7PajAPvVeZjXUcvPrEmdPWryfbg5ZOgw8CBG0bO
5knwfXtcCcm6SBrs6yrFquYcDaZeEI14Ecn+q8cA/+w66Ta7dLQmgwWCFp92kmx5EYphh3NkrXwH
vyB78s2JvIqn7XeuudnzLMKBaqa0UyhVYtThCF0YCjwtH8V5bMy7vMypwcCiy4QC984Runq/M1Pb
a98NdhkH3y+zL8MlkZ3reQGnO+/o2PeKf6y6ukqcdcsH+qwPH9DeLG65QlWK9zXzP8YRDaueRRnT
2wOqDG8J3zJlpSX1WcaqyEM8QyBaP3ZoVURxM1zoDDlFmmtnUDd9xWSJBIWC1Ey1654CgoR2th2S
lQR2MWzsgBmwR4cwzwg7mO5yVAKMW66m4VkUV7t5bk7fEg/FpBsFxf+fYbCnMakZCqtsYCYSz2I2
RfYpH0TFSlzBIGR1dFYES3dj1TT+tqcr88mF6sQ/cXpasiNgKdjabIWwdmEj2TXU6UT/qeQrpUp7
eiEr7LSnqQqrPY7ViIpIec6uNBwYiRnqmjg/VEZFqUEERxqlyGz701Rc0vgIBSdr6sGDdZaM8U3P
e2e3J89SkZIRKIq33Jl4U+2PKIq4vogFa2eOeCZELdu3RevWJzSjs/xar5zubtciw5QJERGHmyQR
L6OJtOwwGFabRNU2Nc2B8/5qwkshoMU5OJcVzde9mzz8/qhWTwJ+6C+FEEqn1OsMWFKxYCvSft77
ZQ6dkGVTtDU9ahpis8+WA9WuzKwAQRpyIM8HtqYKfF5xX+xgI3OSjRaNUcSII7BSIeB+he8ZAgOu
VVVgT+DNfJ+8rgijv+qcCiOMXI2A9UjrZYKYMyozDsvupLXk5quWxzB3i2uUBMVW9fQRrpbPFrQl
xh8Nh8c1cEb/8BMV6/OBsp+yb3bRfBYzSw+uE4KESfWIvjRaZyohmYyGQLSUzPWG8y/s0VFztXXc
/teZxPqffjo68VMrqFRGRN4tOiSlJOwE+GEm6NDqPD6Kid6CbuMHvuUrN4ejPGZygpbGacIX7RdX
PgPwn3uTA2CTWckH2N6tRgkO41j8C7f59czVOYtihFH55H1STqQNWR2vDQn0/AXtogztfNKzrsP6
tGQ8k4X+BX2gZ2aKHGjLcQ4diKMZ00oxavB7ICfjn3fS3okwkA8KqPKGVswRva4fU51y0pabNvNW
K3wmClTOXuGmTjoZ1uKNmmVzhkvsc2hbmTxoRclV+boMkHvFpnQ1fsBaAog6S5KC/6RuVmBYgvWX
rPuXXeHhJ6N/vsyIJVtJBEcb+dAG29hJyw+HIRjnxNYqf9zC+7oJNvQtJhRkeYG+uWZh50FcgEaD
AeTUAurokrg2zwiXpe8dTJs0ah601g1upVUA09pTdNetwqlNDb+RXFtG5bPGm5NyKerxkAPfsZZi
wJ6hQM9fvYTJLbTKDMMpPZngAUv+mlqkui3WoiH/gxXQAmHei3UwIdnQsZ6bCOqni7I7BPMOnDO0
m4JgQ4orx8b4bKQpJDS/I9XCVc9WPsrcKOFVvWTU1bnANmLEhakMpbk2fVzUCdVdrbPyo76TzIgZ
1cKL6VAqfSsUa6oifHpztuZ0wxQOTFS2atc/7fHFTGdvUi4VVu0KEEl8cBeY3Sq0zi4E68oUOxrI
WjKdr5VLsb2rAIbCLYVothmyf0vpIlpiTVQREdUSKL6Kv9Q+EE6i8PnbFj1jkTTfbS9BBVQPKWxI
Qn1BNccqf13mVE836jJ98XNyOLqS9FftqypACZ05FL47C0sssdfClg5atXRRxIJ/Vb0+YTwh5JGx
cslu9OwQDcOBvP+I8Mj9+Q798jBzi76zUFnnr/uCinSHae0uDzYXvpW3WWbRo5/cXo9LIEcCkBeP
WiJyUhPKzkON8OH8fFzQaa6zMYHOXtUve0ayp7VUqA+5k8JDc3FSBApCsi2T1USqvO4+BnlWLQbb
+IsOjdYsiMYfEkl/+y9Ipvfy9ODLAFunp6EnrN9XWYcIhzVCyXeKRySou2+SGKvLdpeGpqV+NclX
smxKJNBtLpjns2GPqPdV/oEnju2A952pvxhXpzXe7GG7/ClSZ2ubu80XrYGAbepxOd/AafjOVRez
dEkNKcmogV4077/EneVLU16NqR8QEMpunPprp4xroPUZ3bp9T67ri/opjRZtnAIpc9dbIcfcBZn4
/1946Uw1NdHs7U5y2eMGBRtMHGKxhWXRlq+YuCxomU+7enqAUInoXtHIq8DUXriqNBWffJ3T9Yfv
/lbEnxjtD9uZa46HKHk6W25akXHv3NRcbmrWhESykXJR3aVPDv/GwJ5yS4/5jUkjO6m1zYtLCG0l
w6Kt9T1UaisMsFa7GjGX08vPoYGcWsQh9CEpO6GRBcTaJPNbQ+X1gzm5hqXqQ3G6UmeQz64mTrQM
e+G9IpAqgiNBpOVwUJCASbheAUfYY9GsFC+5UZwy6qc7fsqkjersyfWS06JF9EdH7VIcrFZc0AO2
WoBl3NgxQCvaPeOmYqcqIe3bIXdsekalT7O+cHvEKixZ2a9I+vr81wTyzjQL3dZddoqJ31DM9WIB
qdZlhiBcTjCi3IyNSFAoS6iuEEM67zjrHSVZRXPKOulPkQhwTZvBEWy2fvhXo7PpDD39VAgEIJgf
/JTXGpmM+Bpt5hy2fGfBSp0TBM8upn2Nq2/yYOkmL0PZKzXLmUXWQt8kwHfi0uRVdzvb8bncS+eM
/AaE8tbYLHjAOWsWoEFLh+WRr0Rm8QeR/R/8waPBJqO1Yd3wgbj/VgX7tJr/L72WnDdqom8edmRZ
ReqcWAKZkhCTg+vXa828TJRti7pq5cpceAXhaW8yOt9NeSnHznezArYWT+wWrd+SUktxMqcr+QaJ
l4cGbpyIwhVZ+jvxcXdVIDXzsKAr+wW062JsnpCw2MLFL4kbLdVqCvjAhxDwISbrG0cKELSTdDpo
00toQnNkrh4Eg8hGT7WDRrEJpAuuhLFM4wJt6J/UrtPjOAlBdQRAiedS2X2iR5GzAN9SmkiqoyuA
P3dJaUwA+t2z/6lHIRt+2cAYOK2wiy+/2MlSlbdkiWPooinmVqbywZYswxWJLJQy4hbWdyQWXATa
smu7UEHEoSokP3jd0ge0IXKqgsdHPLpVyaR7STB+TlOFhCOlToDRbzctihiMtj7DdLE/x/hGZxB6
1DIQOfRemtuuAwkpnJWLbsep3DvaXzQ6fDeXQ3iTPZHe2L6tsj3L0SOCA/Na32ulGuY1D4vywL4G
NRrDJBy9crdRjh+T4Tnc6W1gjVu0pKwU5xIkOFgoV6nYsdmWecYmnZwPshmCKqJgAO0EkThJ4bY1
7v+b33GoT7xJEgrIry87gqQ7XIqlOBn8NZqNoxwI7Hfffas4DZwiRaEgQ6G4D2JAgJPciPlCZOSE
DGIukTGKCumN7WdV+VJuTbpJIsNLvjCJZQ4U0JzcGCifH+PJNYucqV2d3GqUrXYAw/Txag4pZn1o
f+7mm/XH06Vi9X+kD1yEJKckVjPpQLy7C7KMjU1GXSFQZFe8dmhZqmoMPwIeWh4JxDYTfjaDwScB
JlltdxlBUrOtRrh9tUbol1aY1iusHnZRS2iLxRrpd9Yv30vXygIoWrGHkmIYir/AtEZcoUQ+kqP9
+EUJQBWTFxkWdvUqNGpIiOnQA/kJNVjM5t0xZsC7QU6VR5g5c2jz3WeM2/4VAa+hLdFrMWhJnhif
5jo41v8WIgVtEcE+V2qBa/mtrtgm8JkfiWX+CjkaDSFmf8jPiYSO4mztLVzPQNw4oyHd2pi3m0AF
HNWCyZLRACjUNMk8TZFXf6ChA6RFxPb0N4SoGM1KKqW1xzjkMn7+p0m+KIHnHrcPuVl3cL3dCVnS
oaaPcHH3riUdxSJGNYzUAEiN6lgQuAYm70ls2eq68pvlILZ6NnzQDyg7rxJ+Ykdd+mXQ3jZ70lWg
igyqj9srm7bC10EE8VjpCN7+yxGhz6Lk5D2W1R06G/6WWe0cYdsTVMc0SOltVKLNjudcBcPe0izT
u0TzD+KPqElMHQeflQgStZkP1F4yqiKDkmEvRsk0tQpzC5oNfTnrwsmzF9C2a8MLgZIwqIUmK6UP
h96ytA+JMyZwq0uXGqF7vStkr7Hn/56iicntxeFU7FWeiy8eKpnHH25oL5AZMKYtSzumur+/dI/d
zj++JbNhFfn73mj9khOi+Z8pQbJ31zpVMtQsXFruTMoeHkAYIqtL2gRXr4FuRGLCMuJA6SMw107m
MnOjSonGLFvXBEF05PsaHDyCIW968lvnXAG9LGV3eu0N2Z92c1/HAJF3wWXfdc3gbg8Y+fIg1Ds/
IdQm8Um98Xyv7CJAhF/xjRviQpMppy7PsfniTWKS1k0IwaB1UzPBWWNH4aALrpK5FBAcsd2bSp13
gUgLjkJ4lGliRsPGt8ylH81d92w22p4XF/qnO3j8DAhftfHhCi6m1b6N/x6Ux2xiL0HcKcQ7DxBx
f6bVpXXJatLSwxPeq8Z6G/GY8ogdGx3A1aqT45CASi9Wstt+E9nJzceec68McyxEBBKe7Ez43mhE
ZeMPBhRXSPyts37sekgusTtm+B+BVEBaBVFGO3LjexEDg1T1mXDwMCI7aPMVTNs4vgrspaauMm0/
cVJsdXgry5GvIUzdgPdlf4X2p+f0T0rQDFxIVjl58l47Twlamg4FegzovFH6LsGV+99koKGinf28
9kwKVSu5H21CH7dvseOHM4L1ej72tvTQixfth3B207bQljg3ue2nFweElpzY4Y9PNphiTyHkFSwG
+rDkhGfwKqcPI7P3MF2zrGpUS1JXjDDFvrlpXmINU+RkfKxHO/KdzOManDH3WV3AtvK38ku9J9rq
YO8LCpp9MOQeLIi/JGeYgMZPBHGOy1QH+pIYXi5nOYVNtE8S0DehyyUgB9V8lA6sdgbZjBE3q7Od
yENdu0E8BK8GBtkMohUBwpDPza7uGqUcYx+HnvcabUBn5elcubgUMdq4XnJpvrKGaavkZmlxHT0Z
JefAkTSvpbjEa29S5LZL1dIVunOYmU3+UrrtnpDdnmnU0lOoQ6kRQCG2Vy1pqVnb3+TDmSfS9g6W
ut+h5TOm5J2LYEqE6Pl9SVXjUy+qq0yX7GOHbXg4V+6uZma2V/PMSLeG6qggsBfYXBIzQ7upXn7a
ckm0AZ5sRXmnkSgZ8T7/qG9XiMAUQzSt9YB+n/QlszHiCkWoeRIRLmJWRH6INa+Y1bjrYf60/jcr
UWiKuAUPhA9ER0eH0xHVgFrJqrvO/ZAK3QX0uxqzjF+Gg89oX/Fkqamr+hnNZAxEOy2bVShbuVM7
UI7DCCXxeZj77N1+MY3WsDJTjCJtUotxgRqwIL+CkQS9W6GIroplkoOo84/9xTNvYQ6rm9/NDFYO
OwnqkpPToySwDcEBafrFdSz57ZgbOSOod/B7n4Aqyzbw6j7ceT8COs0+wf+d/50U3S1nuerG+y78
y+QMlayuqqUz5Fx9zuLKm5Rvwvh57j126l7SoxDUACHFjgpKlRCtaOq0yeNV5FsJCwPCk+ll2AL6
tk840Vge3mRfU2+HX30LDeEcjDVXWwxu0uQz18pbScKbm2wMk4umqO3w/1Fz7e834/1kq7vySVRF
49JxasiXQVK16gYbgCKWdYm5NizpLvFbdXM833s7o7jWBo9dUeLzz221I+SbA/MVRo4wLlMs8l6O
6XuSQu90ZeG9mez4JRDnRFy0ruKGhP/cEVIoqxdyG230Rxp5cMYWmZB/+FqBwlTg+K2G4mgc/lvu
ONHR3/LdN0s+ws3YWuCoV2kGvxaZmyJJ6/ARGsfXEO2VuDthBaD+pn3SDfxswJ/UONsZeYcbeOIx
WVx7/uWBOZ+4Z8LELfo61USiz9edfizibPJ//FpOWG2boIrp7vc0u3SfH7BvSQRQ7fncOzT1DNIW
0DpVkMZMzF/NFi3ALTlep18G1swixYXBUg34fjXKi8ezzhaAm2Dkfp6VBtjw1DunQNOO8FHzul49
r4XS9lMkRhl8j0pVkJfFTp6E34nQSkWR9E9bstvGWwTsfCWOlLAe0hphEql+0kcpiiEht76PAbzh
67YiUXWgwQsTJMIW6wrxjvJXSXeyQAr+LZl60Glar6cGlF2tAN0r2wmCacczH9njMzflWemigqnh
FgSKdhQl296Ow68XfYKkePHBDtVx2MQpRiyBJvDeiVc8E8/rA/pIsJB7W5xvFAOUuP4DH6Ne4Kzb
nRjYuTwMZKFCXyUZ4pn3dFO+giKX2Y0mLHJd8gJnvPu1L0J/RvOiD9G4FZJ7MKb6FVHC63wEHTNq
MexnmfM0+2S1xgbx5b0bDyjnUTxGv3A5DFNWhZkL28YsvoyGPa4Kr+e7+0w8HTm39QXvt102Eefo
MUBqYL2RdcykANl7iEcqTWp19siAtPDplN5eijdEw1HMmL8l7F4qkmAEKI3J8B2JJ9q72uBq1Kmg
0TV5DV7ueSugga4qUJB4svNkrYTyQc3pZ56RskD/lPMl+xddPabwl5RjT0iT5Cp+mNig+1zbBai5
HNMs4Z6LbG4tj5tOkM+R1xg1KmC+O9TRgSfrxEvRZDv0fVO63ctNmg1OeNhtXSbC++Os+ML5dfr6
3W2Mfu9yceDa7QilJxwZxZva6qSFlpsHOYsulp5STXNLgXzvxGonPrl1W+bGYZ21607Yb7z9FBHV
n4Gsj6l4rSSLnW8IAshLdsjiU9s1Z036UmaGig/cDK7wcRY3hM0k1N6VlSdswTfhTLNIZeYs6sHJ
10VR05mwK1dFOcXRt2SC7lRpwetvz4A/yraBGdL4kO8xfjFP0hwviGHmmbkiT/h33pnbIFLlGiJ8
MJ9WSlHCVa1BiJT/rdQH+9C2moDxj2a5dEl1KpcP+QEdsiJMbJT3IRAq4vwIoad5e7OcLbbOcWuZ
ru9wdQrg9YTZ6EF5JyQX0ItyElzT9HU4iTFAJaB1LHRleFpsLa84Lh8Vdl63Z+gV63u4HkMLns5+
6CsNvDIPyPeApRSEbrZq9nZPgStB59U8F4qVv7wwBEsR0bneVSk4XCG/BgDET7OqLi+Kn33nBjc3
kHwKUyip83E2ds74Vc0NFqS4rPSDnjfJd2RvlcQfE0ZglUypGp3xY0MlR4/EyjjzazvTsvy0b5N6
pgExIGZUsgl3kcpvSjiIhF4+iorQcmHhJuRq3xQrYeOyfst7D7j7hNtLpLCWNxlR5XibUJB0G3al
hw4kbl6vhUnuoqiGe4wktUjJn7kavxi+piMu8fDQ0/+7hSmO9i7bQ159uL/10baqmY0MFTfYk2s1
ls3Zm9HfjmzrXF/z5CES0Qf7go+ndXvGiWwPqsa6Ys+BMSagyA9+E4poPIdW6aqLjPsfce/TU4KG
Q8gWOkYevd0BcZaYsKt8HsdsR9Dp/KyZQ7GSVpC7sKxNfbCLvPGYgPgO2VHEZQRz/P9X1BBPoRDo
hH/Dh4IaZtfzhkZfuWzMWDkwB3OHVm4X1R/JIO/alPo+Jy3+p8zGPDpRvrPRGUfOBnN9rR3s7awN
MjbCufNXmnp/vdMHFpmvQ/9B8qXfCDyQJw2af+hRL7AJPPnrFRszB+Mnc/6LHz3DeLngYpGVoEVh
DbwCqjK/qij8Tb9luLMrJkR1vf67V+PS0IsVYzHbfDaU2t1ZT1s9dHgcHfxWEcnqAGmSU8Ul4ArE
60vl9l14Ko0YG29n0L/yZTBy498h0XSZVKPbhnIZiBqA3uv0gqjQ6D829NKm18qFBBNUt3XEbBIr
SUOFAYMkUlgme/gFfjgEcYh908Jxrntzp8339pIY/pU/SpMQV7YbPNcnPAE+nw5Z4kFQH1arC/is
PvxjEJQh4k/YseP1T74QH2SIya3nPTSp4jMU76hxS773uYRz6OxZ7GyKVZlw0Efq7URIp7KTW/ap
kNx3exwZuC94JEGvSa4YJPu7BVmVzZZ+3bpimnb2K5zd/aPag/ji8uOsdyt1JzEaCywzKu6WjEqL
Pim0dPZaTuS/3yXzSgM3idpYJ5owUReQB2xPRfdcMxO7nlww/Efl07TTxbqOcLF9H76EvsYHa2tF
bGVGz+ehIMYMxz6WCW6lPSM51ZbYpm0rP/Bksm8ApURbo/5GegHsTSGg7i9Ub9E8/tsM64/Moaj0
fn8QRYK0Od5bo+CieqxxEPD019fSyFIbZ5GOEw11AT0tAAKuArGsoPGNq+yIRA8vEWOyMBtHgeP9
eK9Yvqmt6W5emR+xqhGtT1nzw7Hup+po1o5KTrAwz7+DOkW5/KTMrooeeOrPhT1v3xPOD3zUps+W
wOVWW83eKpUqjufl5hGxJ726VcuJNPnIlDUpfjLFYT11fauFyNgoazHhAu7udGzURwyn2XquEwt7
wiJ3Tn+ohc2ny+7dqt7gyXTNvypm9P3CDV7KKcSC05WugH54Y/B3ly586R1r5NoMMVNH9H8EheoI
1HHOh1FTd7pyDgy8VIrpJhdxsUx7fFYnso88XXbgEHpH4DMmwl2aDanOWtzx/rqsPi87mW5oxGaR
kjs8jcfkGEZCUhkUxKctzLDT2NNVU8Mr+M6Tu5Gy+9EKJXbsVLlU5DCl7yc7zaybU59b3AZ3jw0W
q8Ya2PqFlnYYboRBHhvQVnALkBqajKAEGHfsEOqCPxCJDDxd9A0KRGA=
`pragma protect end_protected
