-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
gps19+vvpuzWMBxeEbbR6kdZrR+htMJ1V8JUK55BMULVo2fd+2NO8FJuyckuy5YN
e6m+E2ujWzyN9QARsR3W+s1YFLHpJJU0NBw0OQCggdj3Y6kBcFpeXUONyfe+dhOD
oK6UnfTqFf/eqdX1k8F/DUUpPs7r6rU9dku2kyYlXm4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 7075)

`protect DATA_BLOCK
srTgHtaASN51lahXld4Jx22cB8n6UUEog8m8Lsdd3b8f2r4zr5ElhsRWweLNK23X
TGNtUs8WxVywoMHbXnI74ijxTfVTfDQ5h3uqBs2FhWpl9Z8j75f9TRYPml7qq/v1
FJ4vQYO5PGJZRKo76kzCvWzhDbwk7MNo1i/anLyLrczaB+BkesmkLdK/M48wDbZ9
HWaWUNGQWhdBHu8ax7CkmOkwYyK5FeJycFscACsEno8IeiS4HVvWaWq49K6uYnDW
S58Ym7ekPolqmR592gTH4X6SfDkCKUJ7zaUnIOoAiTWeJhyRUZtf/POABKT08XjX
xu7HF1584BxfCRerH4QdtZ6CRpm9WcRLbji68D9TgX4Yrkjavv8CzlXGq4w7O1OC
kQAt4pwCwQVHtiKCSP6Pvt3FUehxD5DDOKPhBLiZw9OHCX73Q+EwzfoFyzOP98Pm
NezeJdyUryHDBYs1vfhKUF/YYKyqhvDLtxUROeSFFfbx9T34aCGPjpRcv7o6k5Sp
h1r2y/C9Hj1+uWUGnK6L41qb9VorCfisKP6NxVzw/PvMuOzeXSnoV9zDhFgybWV5
GO1auJJ97dNsDHEzUv11T8UeKYmYZxBRMWbg8Uqb6BkkWsv9gLq8jiDSgDsZwVws
coJ9V67kZ3ZM4hhq0g+mJrI4i3dyPaum4ZB9Tgum7Ni71KtACEEl1ZSg8DKmCQVx
8UCU8pGQ+V/S4/ADJ4UEGjfX9nmMHWdwg2OzEaRh+Hlcyyr0k/KjciETjKKTVFzw
Wn/1XIPViHwXRZymih8ZQIqWC/Sp/so3vdKEY+eW9xyvaWOSuvt1baAdzkfRg7dI
FcGIa9acFFJjrUVFEXPtCs8yvA7DHKUXvbO/Dr0mu1EHD7YL4gFjXZeQqdN5W6PM
+21vQLmOAIZuH69qXIXNWjjND4A6FoursP+y4+zKWcFqdo3+AOvb5BOzoQBkwlqe
DiDcxs1iu4FzcuyomKYk4dwEEMHrzCxR/2/wMXcdSEmLc4LrLRpG1ko2h/S4otrX
sDIhru3TH6ekwhvn1IuJZmii5UpwBbu/oqAqBQZSm+Eevf29+YRR75nhIPJkdNF8
CaRJasxznuPVUUsUNtAQFa6K0FgZNBERjxCFA0351fJ9poL/+tCZATElWmhgqoTX
Ta8VywSiGGXHvoAW6OW+7c8JQUz1f9klI06BeFqpRq/AP2crzXQQ9empGS2d1fsE
i/BnttWoEo4X1YmehgTN3jgHK3INvqC/2X6IqX9nVI1ksKOpBxHA3OkJdQwHukjh
Rg/PpWx2hVGFzY3K13SgUG77LFnSS9EFH7/FQqBgRtbJ0xuRbG/6fnvPlvBWQmLy
1o5qWIJKGqcLWufpNhMJm8Gml24KA3kl73UH/fmULlO4NX2RXF6DGLYRDZGN2pIC
g7Ch2PdZvhAytjoHD+f4tqwVFRewR+6TPqKeSwVHgVfQcdbUQlDCEiuMUTz/+Sqm
jiCcwzIOFcAIRQWcQHYDZE90h+KuNOlFEviI4GLKH2PAnB0bddFOVlxLDBhxLd2R
CKMXs7Ay1cRNcTZSzvMfBIIY5EOOrjnZorJKdzlg3LU9Gpj724uvekuZCr8q6aZY
Ac4TJJOBhcMVqZoTAg9NlCu5xEMWYbGoXwe+r43Lt4IvV1L7UX4ujHVSwtSMHKRV
fFfUrme06hZiwQKCq0V4xU/B6cF9SswGNf6NVH3P8iuspDMWk38/hmf2CiD/RO6h
Zxdr92e3amyJ2oE2uxOEwY9yMXw7ONabFRzteXjYNS0nJmNCNY0RdWw6CygIdGIR
Bfk8JYMUJ/FWCHfNYRJPS709qgKnnb6SRNCBqByEJSr5RFL70gfdtTLFCayIqHyg
ofCeQB74v/M6TSrCfqIw+v5bCEzuW5QZgEoAz4DBqyBY7N8VPeoilslY3ADsGcPa
9IPC034Kbz036+bxcpuRWHc8tkQ7uKlY2bbFk8lmDA0NpI/XEWk2Omx1IQcem/0s
iDJDuNKkgo/jVy3uPjmFeyq/0i7zQqFw9xLCYdJC2swOSeelLBx2Wa7ssYpRRhHk
259Rv+A8ZlvJ9fjP0rEGWIlwI3GN39MOfZPUHc5r6foYoImY93xy3s/vrJDwA8nL
Ha0XUip5hcjmAeK/nszVVjoBGJUQAXGAyunobJFBKddqgu51+Uf+NGsswEuxHaD+
aPgorPg/uKopu880f580cdKCckl5bgT2a4yvngvF6VQF14Ti78AT6Rzfiseh+el3
vFLNGmilLcKu1UOmAy7t0Ngyjxu5uxzhiejN6Ntisi6gAt1HshC0OVIbxsZNLA6l
JF5WP26OzT3K0aUl2p9iXzhOVg2ffyaHkUk7bONLx6Q0daJvRH+6F4OnzsDoBXq5
Su22fZfRiB59kKJXKP70qJkbrdD939QVXu9kQ49oSaCeSLDRh8YLXd9f1yk1n2gJ
MEWi0Te/KScxrJbIBCKBeklN1ArrfULH8r81vOgHPC4zV87PvH3oesIGFu6rpc8+
NgD+nFlAf5mhL32eDkEz3AWU2qH0plUBzS2C5Sg2DQ2TAHSLsKs+8IX4thh9Nqi6
3pErrkWHOFtIiQWZe8HI4WtgnCnR+lMJgYeaZzYkoIRR2OJv9h9A9gb2hasIxfsM
skKLiTU3sOGoN48/9FkR4PnqxS2rTycwy1c6UywcoWQR9siOct4KR2m3jhkFZ1tW
5YR0iVUZ9KN3XZME9XJw4OW9CDyIMQht3cluTWMCx1bFUazJcxHRu/B5XT8/yaFs
r+Ex6v5ZI9QIQwvNTQ+cl8XUNQUR0XOUF98Tu+tkdES6knoLk9FKc24k5utIi231
BhAfBfL7jpVcVP56S4ujXuAx0iORPzwKNVM0X5rIlXt6MSTr1O3uWYNc2etETClA
ngXfhx/wyz54qGGqOV1NxmN1vUbFSBB8OPnV4CKMuIAvMfwlewfT5ksWjZsj3N/s
dQj4ysdVTANo3b/Tq6/A0Fa5cn8Kz3lGaCvvJz0zVfSPRsNc1sL6uTryAvgnkM5N
5VpTuHO+/SXXs1AOuvlZFi1cFk8jsYIYAOR+7aGLvncmrAl5R0W+hPgU9urPatuI
PA264R0uxXYagaNQIDH/0DT8R8rN7N/HNajHi7M4XVPLRxVGfr4Gn3dqjeyAzTWu
aHYEBwqeGigMD7VHPdRIFbi8aziGxZb5UWQVcXOIJXBpHs/+fE7yLR4DFej0EIhf
CTI00DrKXeNZ1z4w0uJFOvingZBM91upKHLg+yqaLPZiLKf9eEsLSr+oSSRhkQPq
VbNR9bDJzTZQzVZ6oXULGOj4sa/umBuGKPLYBfH7y2ChJ8InXkKW8p1gN2uYajm7
a/2HUiuvt/9IDX5niqYgKNVPkAgGSzNAsswQgjnBB6wc1TmwWHvrV/uCspb5cfyg
hLcnLPkxYwcXZqISdKbnVrcv1NndYtLTltUTByBY7WSXaPtDHJaIPqvO4xwVo+T3
vPi43dQmWLTPuQN3ILRWMJVpBcgOdqL93OensUvzyEFCW4julhL/u2r6i/UETRtB
SYBYGolic1qTI7TJ8eoG0uIvTwdKEa2PxaDROTYgIn+hqy2tH4OApJi9kjNKEKTK
iJxUtrJuQiXx0foxi2l00YqVirU5a45MOYNGqGaGu5ta3nJ03DUvtNOFwWOIky6P
wubgxcjsOkfArsLJihYxdGCxkAqSjFoZv5wZpvclaF4ib64JtGdyQvY0vdtKHmJe
Qk5ioOwwRzHiE22JeYix2jb/hhNoeqeIbeMoFasZLQ4VlVOERQ/hkJyjW8lWJ2UJ
wrLKP302dwvnLOraxipl/d7Z4tGGvYezsJpy7TQwrXo5wGKd31L/0js5RlH1tjXx
8746QW4br1AXP1AKSWCQoS1n3pPvPHhLbPsdopgltj+u/2IO8eDrl1KqXaK7SaOY
WrdWCh2z6qjxO8FfDdqoTYrvxc2/2zI6CKbK5MuRCY7qdNphkBJoG822Avf/YN7B
yKtZNBiN2YIMbLkz/dOLF9LfN5vvGyNJNJUOpBPxrvk6fQAPVnHVMDjC+T5VAGF4
VUsgzRb88n3GjbapTDCRSLAek5by3veAjhjU1UPbrA4vCGwtDshjITLYoHbqk2qO
OFw3YzrKdENmoBsnApb7ddEYj4d2WOwtLE8lMYlatadAJOQIN4jE5bWBgOqV/Go7
yb5kdgW/L4jJrU/LrhoiPtuyS7TJoMprHfgO1yBwrUHez9lTiagfoSSlwdYZ0ZEt
DC/t+CpPCgGlw1lMTqMziZEN5toWtd7BtUbgHDadmlG1bv1s1nJbNNUHkYtV0Ah1
sdVHN33E/TGf7LW92MrGCRPoNvxbZjMeShfCbOdDi1yZBC/pNy+F7ibOTysN5G46
fLGGr+XDxJN6LEk7gNjgMl7d3ClLsRjWLoJFs+0lCDslKK/xwoCB4IC0L7EXzvOi
pi/mvjl/nueOtEzcJVStqQZjH2ub3/Gqf9OuTgG50VJTfJaB8GpXYMhk8Uttbs0y
L20xKp+KGRMdya23ihaUkrXq7XWQyFin66DcHW0o4wZ1C4LvXPlxwD7f45uXJHyb
WoNB+uoj6+yFcUcucGaF6u2rNtlHTzr6KcY8+6LBKchQw05h8fq4Q7dOnFwE1A2J
2iPoR/d1qQ9mxspDxxCo5RgMTT7A5okaIB6x3YM5saLrFVMfRS+sAZ8NWrhrHFEA
MYofPl4OwMZS9/9MiovKGG/L+7JGaUlY9pWV+bZP+j1iw6WY/cI4uzQh111v8//3
GEKRlXGk74qQCvD4zZNre4JGKUCiyXurmJdDKcAOxdpgBR3AqRjf+n2NBGSMuoaf
hFyhRhlkqsnCEPPzabdxY4jMn8Z47pDUNE9FfMjHwak/vNmMOjFsQlOjdtx5IA2C
HD/tmdwbcSl6lmdMFK1V55DtblqxhmcAn+iCYI9G6WAWj/zKWgot2tK7XaWod0TV
W9qKzXQouxm/01rAWhtqR6s5GbUwxevZ98jrB7IuxWF3m7+OSeFvd/KOaOGSeshS
Ry88XClUVty5ZKXrvMBix95Sx1qGo+jZ2ZLO+DI18M8QyfdsqLeAa9hxcR9yL/JG
auq8LHPYdfc/rHH9AGm9/PvwKGQ18Kn3Q6IfjjHQ6VdNO6KEeD2+492wlmJhKrxi
HuGDHjqdW+nDzh6yInAU/XmaMa0ge/o0tvvvGT37CGTUU3HPKK2sgiue38qHF/yL
brNG4SVkZ6iiOupJrUeys/rJrjM17VjkOxu2CPV/6HQ0+s5r/HtJK89pBBjQHpvt
TSykdge41yAaS23ZqCqCU628PBGtUQUJIyQrnhSrrjjYFT8l8Ep6S6IZFopC4Qq5
qA0A43OfWMmPXZ/1ylM+mNO2QbwTl05SN1CXtEYLf6v3cfWbcdIc0QbHspnmkDj+
1BF9JT0N53LiFQL9ew9pMtz/wSIQDJJPgw1DAZ2u0fciDd6CfGmCrVnjaSCbIUI6
HMwUCvOtKOUoxS3uU9Kw6rjTLAt4Fwo4ytryDfCIaASHH9dGEGebSmpl+nrZbBtT
Om9Rvd6Xk/60fiUzKjdn+GmVZhtSFyeimiFwmERe1cILrZX/F8OoEEizoL93aRxj
2T9wuBujCGjZ4LUgO4kdYFCbUamA9ZUxH/bhVVGL2FoDyGsF5uwBh0AwwSsUx16Y
5mCNTen2pfoDJUZnEstZjGKjYdJ7LqPnR1jSCRCV1ZWVAkcq72rvHoyDX/ZNR8Op
o4txdEVW4jzBtcdXWxvO5tJfB1m17B7bYLabthc2aOn/hqMrN+XfACZO/cR24zpz
+jQ1xlUYaUmkAkFsSkeiyq4yh6/3jCp0I6/4j6mzs1EGRJuMMyhqwJ0TsbM8c89Y
TqjtU1a/CymsPJcCf17Z8+20nckbV3xBqy6A//uBvthMzMXimdnmUiPDIXDwBvSU
JCz8Ykm5SLCw8O1vtGxJP63K7en/y1cNUj2yReeLoH2T4uGDInAkfu9zSCihfymE
/1Z5CQzh8/cHO+jpX5t1NYcbkfJGFLNHXQyLeVmWSGG0wIwRIEOrsElSG+VojIko
2R2zHfUFvE8Dl1PwnyDalMTYwWXeC9pZe0nr90b7SsBkyA7M6ngm2Ov91eEpcMpF
Gg/36o6oW9WaZ/DMJGR0YXmSDDhytjxcdbepSKRIoOADuWIx45uI38R3KvZLLFJs
Zi/mu2I4F5UnTXBR94nIoOz8IFHxOczhQh8NiPCXPi6CP9Jtf9AtLute78/QgEJI
D8MkRtdA3UDnxgKDNaNwhvV2jxVoxWiwRC7qlahKhZ3rFK6ZnIYfv0FzqmUhyGQz
DVJ66EE2d/uY+lwB6xAgPsZhrPvYqJhpz3V0qiSK0MW8ITKDV2AU7X8DAxfffJ0b
DFoohdDwuL2ObFlFXzkaITZBOMTSQEsAAm4gKwUoEosurjGLn8hXI3Upt0FgNTH7
1iYTj+2Ix/VII25+2M7fiHL3TwshV5kHDa3G6uXHSn14237/KB7GZH8JKcH8sAdW
mfnPjj/qIj7OLl5uvGL53V2Zc9JY6Fdeqw4/FP9wZy4Me4MOs7KCEixpzsCexOfO
m/74oqRk736UV5iwGnr00qH/MTntHrBg6QKTURZB3gmd5PMYgIl5AyuyD+Q+omKA
/pg5izFYwlParexfKwRUY3Jwa7L6TtML6DEcnrnGwOXYuRyxKI5VPfLHW8h/17ur
WMGi3btOYEj590V51gUyWeS1pckKYJUdf86/dQGlAMNdrhbz2eQwYpRR6g7trmvq
o69P6+nu8xySaWlrXNJYU6ULlOOu1T4PuFTH6N97KdZt8sBV087vvcaxAJsQfMwK
5S+hTOrH97LGlrQmBPjgkwsEIZ1Pkidb0kUVAKQ7F0Snz9FaFxuwp32zgtM1gnB5
gv5zvZd9BGumW1R2Ha363+mxaqd+j5sghHv6dhmfE2r1IhWodO28e0C0oi8u9/ZA
IO1TbfsKKzq56uyG6FzjclXIJIj0Rw9AbSMaCZGsKGLQr0OCsGrdWxnL546FPZMq
tphEL7+Ad6pHiAgmBvV1ITXNhZ81EAEXBAqdcnKu77QOUG7vBkDTQmHXWRBUJvku
AdAvtmF8a8qXbR1BpBcmNTFmL0+HyCEc9Yly0L6t0yPtNI+6r5VyZBO210oTTfEq
XWgJD7qav17JZ3lc6smVJkrem4KUZQT4dtoMsLuVo0hBg8V0W/8WiWve5nLFsjy6
aG/GHkrXkrOKEE6zg8wzwvM3073qN1t0wVw/DFvGUN76MHMoucitTNJry9y49/L5
65Qk3IdMwRp1wpyJ8vsSn7uHFEeP5HV5gcw8zhSO1Pt48NQg09fRq9bqwbxudZc7
d9ENexWclPRvb9EsttiD4TzJ0/TLQ9GSEAVT7kekb4fq7PWycnRM/Gc6QPTTFBj0
4ZwhzX9O0IcQgwRWHeBUDZCWUG1cODYAGvxaqInkfdRqtuCO4iTMgNqfpUkheAMI
pKHdBXfGQDcsQOEeMjydiYUXzy3dEYIYeW0SZZ2PA0klZcqd85Iqg7PfSwjnnG/d
nA4NrbF42vxEHyctV4AFpIefK20t37bfx/V0zS1hzcSuDDVuJldpgS3wI/doJYF3
6m5g+6jYuz7Y/NPNajD4LR690B+nXJPD+9DQ5lmAumn7/HtBT2/Uqhs5a1Yec45S
NvOW6R/BfSly/tl92sRulFq/xG6juMBUCz4XYPRToBPUdBBWQMIsyUtkkuABw/Tj
4UYS1sZcR9LoZc3xZvJoyOMIe9tStISpJwwHsXjClyQ5JjlEsdh37yBntSAheUiI
JGmln1hgWIrJc583fVy8OUyQ/koCNeR3KPIzJgifIkruGjZXn4oULswMwVC6mhB7
cqTmCovkBfBOk0I+qY/ZzsoHi3/zReZ4fqlAEKGaoh6RqOAKWXHzyZRKtGWJ7Scm
DefnvAK1owclJrA9oGg48uvwL/gR0T65slj18EGpIozYwibJ18JNqjk55HZnU0GA
TNVDbIEogMNZihlL5H5dyrWkHLX9WTmzUVkGJOlwdsBoPtdOvVLpu4I2r1cbEgFG
pll7FWvJnAG22fXDJDppNMYe5SwNIA+3pM41QKasLBbjusO/F7+Or4IlwTg/Lgij
CSAz+7nURKK0hoyWX2ralVYVnY2oACE/0BR7g3EOa8LbTTa8LdcTzN+FvzYJ7uJW
6zImc5+XK6JWw5mIl+qRzf8KZQNKbZsnJsKZRS8apo1G+GqQI0q2swIFeXdSLcXp
+0oCMZJFk/U8dM6i+Um/EkXtqs0g5dpiFDp8YpRvs+C1agfshxzgRZ5E0mPXP+ij
X9/OVNxMKL3j0ragErOvO8NBi9KaqDsQIlePby8R7D6l4Nxf3f+lFLqCJAGvUe4A
Br5Oo4Pw9vILOaQ3alPESe7c/B1KqIYFE9NViAm/6o7WGBBuOfkdvc3dbYlHaVRj
8DPzsZP05824O8pCiNdzYpVU/IiOmkNifT/7arJILG0Ya8C6qEXJPGNXCNQRSjgE
eEuEiBhkYQQph36cMGTs0HSUCk7+jHNgxuidCRYhd5xzKwoVC8AM5UqWvuKqz5tM
IaEzb+ajuS/U1wRlKKOAdyHSdIt7sbGaxly9KDXbfv8IsMl2xKy+orh3ud1UT6OQ
vpkT0lx1Md+GdQZ6i8L75QvpVOBDtF8pek27PjLMbsBYlxcljR8DtzxyMtY1DwRC
ahZw0Boa3uYzOZR03r2eYzJ6tyh5FdXgdRFSQMy5f+JclBpsGD2xw/AASSKxYwtu
nMTuw44fbXjfYhDYsypRfy4qakbR/XV3h7k1Ryh1CFg8Lmm+8WDLI33eE9GVOQJU
k79KXs6VmpERTg5JdCE1ZkZWlPW95jPtA2tGnhJCSgmOsf+PKvtp2kexDM7qAd4w
yTveun09urrqRY4XrL7xuuV5hopKi4LaCXBAOPqFCMY31FbRL8MrZcAxVycs83O/
zyBRwR64VOZJHag2rdR28uj/5g5hL0xALb2yhKNjC9eA4BYJZPdoi5EmmZtwThlp
IiWk6TjVm2mTFh8CgeP34vw3byLr5zmM6bZraXha8eLdM5oloqV18CFZMmhURrsK
APjItEwdLspodOH3+dFSFbJkECYI1hpDXEbA2n2a1sdtS43PcbPF5pE+1xwqboQd
b2hrmP2AbQq1AqTmiBbd2k6bjqQ6EAomxVz29m4hpg1F5jSUoFxj8A04JkU319vE
TeNiVM5MPzV053BbB8bOHC483qBUuVYUIb0/8r66vFH3VynbbnYeuRm2dvU5SOKY
ZmLm/x8S09B2lspFR/OTAkW/VR9qbDqzJnEJwm9x4bsntXi4j55wBTnBpSjCDIGE
PMEKKThwpCJ01pgg4pwrh1Vueue2XC2UpWKfOg/VmXDpRr0BshyBpSPQ/16A0dmj
HXkH0x+T3kwRkZ8t3sf/ATO8fadt2KuAKHYaSaypVGpZrJPSDYCABCiX+eizFVpY
J8HeuYOvbuA+k/zl8JO89z8ntkOn4SszoCuxzy8I3w8/LQX+suitG3J08t1Bxrgf
`protect END_PROTECTED