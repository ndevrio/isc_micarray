// cic.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module cic (
		input  wire [1:0]  in_error,          //  av_st_in.error
		input  wire        in_valid,          //          .valid
		output wire        in_ready,          //          .ready
		input  wire [0:0]  in0_data,          //          .in0_data
		input  wire [0:0]  in1_data,          //          .in1_data
		input  wire [0:0]  in2_data,          //          .in2_data
		input  wire [0:0]  in3_data,          //          .in3_data
		input  wire [0:0]  in4_data,          //          .in4_data
		input  wire [0:0]  in5_data,          //          .in5_data
		input  wire [0:0]  in6_data,          //          .in6_data
		input  wire [0:0]  in7_data,          //          .in7_data
		input  wire [0:0]  in8_data,          //          .in8_data
		output wire [18:0] out_data,          // av_st_out.out_data
		output wire [1:0]  out_error,         //          .error
		output wire        out_valid,         //          .valid
		input  wire        out_ready,         //          .ready
		output wire        out_startofpacket, //          .startofpacket
		output wire        out_endofpacket,   //          .endofpacket
		output wire [3:0]  out_channel,       //          .channel
		input  wire        clk,               //     clock.clk
		input  wire        reset_n            //     reset.reset_n
	);

	cic_cic_ii_0 cic_ii_0 (
		.clk               (clk),               //     clock.clk
		.reset_n           (reset_n),           //     reset.reset_n
		.in_error          (in_error),          //  av_st_in.error
		.in_valid          (in_valid),          //          .valid
		.in_ready          (in_ready),          //          .ready
		.in0_data          (in0_data),          //          .in0_data
		.in1_data          (in1_data),          //          .in1_data
		.in2_data          (in2_data),          //          .in2_data
		.in3_data          (in3_data),          //          .in3_data
		.in4_data          (in4_data),          //          .in4_data
		.in5_data          (in5_data),          //          .in5_data
		.in6_data          (in6_data),          //          .in6_data
		.in7_data          (in7_data),          //          .in7_data
		.in8_data          (in8_data),          //          .in8_data
		.out_data          (out_data),          // av_st_out.out_data
		.out_error         (out_error),         //          .error
		.out_valid         (out_valid),         //          .valid
		.out_ready         (out_ready),         //          .ready
		.out_startofpacket (out_startofpacket), //          .startofpacket
		.out_endofpacket   (out_endofpacket),   //          .endofpacket
		.out_channel       (out_channel),       //          .channel
		.clken             (1'b1)               // (terminated)
	);

endmodule
