// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H)3+NS9[HW-G\?U_!\G+PY49MVJ]1<,(B4KVG =)K QE/H, [WZ9PQ@  
H_LE8L$%@;4@?B%'\#(ER(/_EBQV^EN;F9$+ZQ,<M21-GDA%83BX0I0  
H=:.RF\TNW(;1-7H@!I33-?>[LV=X49ZR#W%3[M:?#I"JM\E[,;!U@0  
H19CB]N9]6 CU&7Q%3GB);+&AR35"F@]RS)5.Z&&L-/-6(E#&XNP[RP  
H3&JJHP ,)/_+)!Z8A;%*5F;D)P\>\62IF]]60[*S6:ZM,_/482M>JP  
`pragma protect encoding=(enctype="uuencode",bytes=672         )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@ST6X$\.?JJ_\$^BI&8,(T8\?PK$\QGZ&)=KX%+.WB4X 
@9Y6$D!7*"Y8*R(YD.--DQB]R%:N ]'W8FCMP4V!B^,$ 
@U" B_9.HLAX#,NT1HPJV>L7B"P[-U$<!=RB 4A"PCP8 
@+6[?0TQ?,K6B90\4BG%=,:#?9.*GG8N90Y\79]1UGS( 
@'),J&P<'Y#?S]/R,ED08?*=!-GOTR1 (B$VSNI>3]LL 
@5<(V<W1@-SU72*?^/E,!^0Z8;TTJ.2:@UN"AM7S(@E8 
@G)Q/&0<::3B0G:5Y*D]GW6SQ3^%(7B.H1)U.'H]X=EL 
@Z1T6>(-7D$-4MZ/>030UB&<<&3&L%53M%)U:()822]< 
@0 = !/XA_Y]@4^@7_'X<^H=#NT%]>XCW<67KGG:47;, 
@=59GSHYK;S"#6I^YCG\'P G%'I-()IP[+-)[!L3QYW\ 
@JGK5;^7=;.0AL%*C^S14=/R!IRAY+@E'\]U'?^!U6$D 
@GD#D/=X Z[[89;<X_W0_LW\D+C&9;)L\%2B#08^T0V< 
@E5*"V7&J@>84#N8JY5\J]YWWX8,,R</=J.D7=A(NG_D 
@FBIQUIOW6OV=3;<Q41!TE=,0OW;<D:H[U"BXN8>[Q:\ 
@B> _>D:WS8'S<?_-$?O^)C)2 R&HYQ]#M9N8LD=/NC  
@\17^-MDO]\Y+\:0.:!O2E>\T4U+W##1)L;:Q_/[XI"4 
@\N;2;7WW4987OX[@1%E*]71'5J"<[7;F+!<WB/X4TVX 
@&R:<>*VAG37(A$:W7V&C0?Y*522?Q4E6Z0];+5Q,$*L 
@"G3J6P(#>$[WE*V&S5_XJ:B;QX 24@7TNS,#"@[]"G\ 
@;89(P;SQF:J]BKH24\=G#(Y+"]B^O>VGKH-RL0/Y "< 
0I?FPXN5Q#I/X9^2)L#*6IP  
0O)DE]^V*F)*.[K8"H(;_B0  
`pragma protect end_protected
