// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Ddp9vDvRlKJ9QvYJXhcSCEyIXSNuNCKootVWTKVvoaFhVxbYJZsK4D7ExbeKc5l3tKK6rDgmFFwp
XUERgMN1WLTkYgaAMYHs1K8tEYlpaVxol9Pv4gYr1gVLNOGZXUFjEcUWqO8cryfa2yWF0LF7XSKO
oqu/Hgcxk/NxDg1c3KzA8iitNIOmav4jFslCm6jWuU8SBP/vj9/R7vnQHHF4FDil8L4gI8cXYLbo
m9rN82uYkMDh2Ap0QIYZJxEIB7u7qrie+1BYknt21K/LWCfpKSGTkCXK8GuC49AXLg372eqBuYpm
1/UYnS0kOXW28QruAp25ceYGlT/OF6oluXpMtw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 2912)
b73J+hCsq04ivcnmuKj5DkewVk9n8HUE60XlDvZ4anOj7G1eoii5Kvxg0gkkCcbk/NFOfHrdslgb
YQgNbfpQhSnf2S36Ym3k/dNl9/bGXkoI3jADPk14Uc4kXhpNTmWJ+Unsvb4oaUCprET4C69UOYj9
PBDz5QSBjYqUJRx6Gt/z0g37vGdrE2FvFbmtP7tmJ4l0vOko8X3A9sS3LedioQSRSSLNvbU3qlhP
6co3qCG479NIS0qWo5p08ZpTCXQ7yUy8/YSy08u4un/Whdq4I0snC4vFTKQoSgj+UBjksN9MXYJK
wc32PVl+TZlBc7SM0tXzXD1JxmPQP6TU7EcSkuPgpo7E6xQjBZzuu7Ey/Ysxo0At60ZvrHg9aw7B
p4G7+9UAPhulGmB8SHv5my8oxCWvMmjlYqJ41KlLrtw/9AfIjTO8dZnH0Q5r40277xMTZIBGnrOi
tygiPSz30cFIuolUB1q8Q3jupkXu068RNEh904t0s995gqNiQTS4JScrECHIilSWSe2ic1K8KM60
9NE0R/W/vWbYz1A/t/Rw9rUjE1Dp0vkHrrcPCI4I9rykiQiMa2eL5Km5YCVOb9/iDzwvKHZEYmqM
mV6rkgioNuoa/SYVO3p6MLt4qdEBxtT0g8CdmKMKyCILg4c5fdorWPHc8ozU6ObFngUownEthGek
dZAxSvHIACeNSvp2DtyZQrg+XoARLm5Cj/DDGx/oGeVO4P1LZxkNLIGeGch0sz9KNNYD82ahE0S7
nwyaLcvSsmtKFuGo9Fp9ljWQA5OOR7Gm8Mzc8xuavRfRDLQW48CpwZqYA+ECtAmiNVzehz/Ck/rl
VpVukdU0SKZiN55gokc9AJJl08KV2gZNgsPuGaP1flrzPG0X98VpTsw0HIwHT2QZnLpUxKvKqdS1
uU6dJyTvJU7pp8B5YhLyxkgTIIg1sFQg77IrrXKv0VwI0i3cfqX70IujSFvIdhh5Lffhw4M/snDF
WOxwpDZBXRzGpeoaxoBHz4yo1qGx8riJDoTg2RxpUCvV3X0M8eNNiFJEFPChcXvkY8NOoRkQfJj8
9L3oJXXEjIIA6eK3zt6AVB59nkn5yp+1GwDCd0DLSqD4LxRVluzUHOGGmZrsX2VTbzE5nOTQI6S9
XsYzX5O40oH07MkmFa8XvYwdSHnRF3SddD6/o+WgKtbqecdkuIJgD/oUj8UH0EOMYWLU5xEltq6u
h04FmRW42/Wb0sckA0nXZL1S8WyLOEXA1QTJ3fF+vrnQoT8QmtoB48Xeqws6dCBmaA4F96ZdoCku
mZZmywqZCJkGwDenuQALkSH3S2HPC9za9KwnPwWbxgIHHsE4DvQIulB/4Q4gCpYbnBoc7m6RhBYp
1Rv7b8uBO8zt0w4f+fcy4IhmFiVUxpNVoK6xbtJQibkV4YbVxB7uVo2RU5kUZ/Hr3VlMviOl8TTo
xTMK3saNtUJeVv6da6a6/TCO3p2Z+Wa4F/XO/arkdT4GkRP1/nnfwXipFKhtprXgJQ7aiVMVnFKy
hTNGjkU4uTf12e3e6Ex/Nmx/5RsJdPc3/gZYLrp5chNLGR3LqYVEMQJlKjczxzlKaqZFIdhKghQi
Nupi/4cN5MM5RZoMDNMbbME1VmvsQvf17vzV0aCjpV4sjm4mwAPI3xqAApHye4sXdUGC+6ZfeVqM
49LbYNEb14t+9y4JKTQLM9oDDf6uhT+r+opVj7huA59oRVi6+qA8aMGyD+Pq9XHWbKoawHuXBFFb
AGNtQ7TS5/iMPz7XiYV0+Wts0SVJf7uFsWcuQT2dyKsDqq+GlhBh85zNdqFJQuVUh2UUitYO+sVr
d3jVbSzCN57bmbrGD9446gHhN0jdfImxs2cquXaKyQUAktTx2+2QGyioWXx5ztAeTAMHdaJ9eRRv
SlQAlsBxTYvHFrv5xxs0gtPt8pMKy9zdclPUzDlB/fIxQwfoQjmxyO5d5f12UBspreoNtIDqS2Ek
dnF/w7NB7TMAzp7xbHxf7OWryFgOGSbYzc4bEWM2TzekazW5zonHQP5nNghx9co5QjTxeaeZwnfL
J3yT3bpI6MvN9MOPezY9SOzDeCp0Tw01QKtUrU46vIJlmSBg1yaNh2lo01xoyPdErkH4oM0pn0ZY
iMF2yCLbfrEqmZrLQWVk+1mlXEUjWyWymVk3AOzVNlwlcNZWKtaV5UfJp5IOnXl/Yx7EuDGtMC6H
1YxA9mwjMsfOBqwNgEzN9dKZFAj/deimS9E1Ps+3Ilx7/ACpZfLRxlRoDVDQWAgaHxydXFDtCrKB
pqQvH2PRaOTUt3dWrk4I5poRFK/MlKoloHNP7hoo/jd68Ble0bl/6sIJDbru5662va4ujT7gTUmn
RVrFnrpas/BBuZV/aNoC3kSwhtgC+41sVszfdRgR0DC3Pq3Y9hDo5ELFXW43GdweSuzTQcPQ4A4Q
SpkgEe4LOk99uIMEI/ZBv17NmffCZ6gNSCpFz8r/RQK+qC/aTQSXA13FdRF6BEBFvCMdEAABoOHv
6NlE81dE9rqHVnvGpJzlQAmv8ANGti6iL5g+1OJZ51WagVIT37ZWaavRa0e3tmR9uu6TavbkJd+T
KAZWmSx/jI5eGucHL34BotASvt/vKrYRFboikUXeCpvN1FtpLTCBbpjIckH7bU3J57s1KLDytKmP
bEWdzPrcueezpoFh7V8TGo3zNGQqHXTco1b7QPHskJIXwycwp/g3g1UBsGZooaQEC4vdG35ShebL
t8iB1STZ6N7bCTQG47KVRpzTJ9V6lEHgedHB6gqG3rrkvFxNfULHd5T2b60lanx6TNu0HMhLscaD
n9PGGhojIB19ChEu6bFqwUGD/1ni9sRwFTHJrLxykqYnfpMc0eYesW1fbVXXF8nKPGHp+OdaKCTC
DZKPVOFo2+BBSrJ5VjZJV8b81jN8IZFpnmmdbKa8I7rX4L9CgnkJuBdC/21Cxs1FqCEGZvqI3uAC
Ie6TTRmLfG7C39RWOR87V0hXhSWb0NJmhhqXAhHO2cE42wtlZcf7Om7FkqOyZCg8CUmVcKsWlmyR
mncQfuJzcwZgaItQCbizY7NwM6Jl5rJIgKrqK9cTyzyPEdkLuFcIP4Bz+o23lgnsiSb3OXmhqPms
meUNGfGS91i4U//TVIyZ+0eT7fM9NiQ1r52UL5HQrdxBU0hKzEpX+ZkOk+1ec4jRQ8dM9Soh51+E
zcKrkOHPziq9GWdL7PLo5Addq5xugNvIdL/DUXihOCP2DwCH8ZoEJCp+TgNKHSb4AF4TSTswQa6t
ZwccChOKJaSgG183cNDXyT44kxZs7ewuCx9uwg4IKuVRV8VDpGW22tcSssWxkoD7i3cVYf+FVbSs
GbQuFsKibT+uUQ/e8mTVfZ6aycouapJ7puVhvDtoODBt6sF4zj0OD1BaqLLqY8FYPJa3qAyZAjYS
znwr5p+3h+d/W2fwtxEr55ZXZwiMn84Kv/BWs/mAlIL4wlR7uwxtZARioRTielDd6OOqWnhMK93N
kqNFov6QI9RmNr+8i3ZJBfVDFa2ULo1d3XvzNUBTdj4URpfzTURiuJdEGRyb7Rq4zRKO+JaRZWmA
gXN0oO9fF651mUxi6IE6u8fZ7eEqXdtFeRqZjv6MHEu8UzSMBjvANQwoaiPlVGAr2mIIUVOsvo/d
GlSUIyFA+EYMDKW1BRC1gRxK3MFF0wPYt2w7DMnBvO17tQIT9DRWhTW3Cm8+/mPuNxRZkaTueFhv
/BINfuCvynNOzTdhKrCIXQqnC8nUem1SHT6HioOEKMIolA/QrSvq4lJmFkdTsbIHlYcq08uBh1qu
XUbzFwVOdVd5f7z/gBdFzCissNt/WWS40Jfw+Ikeq2gadGMCMKbVD5PlQZtu8VZuHLGx4hGXqc9X
WXRG4a8=
`pragma protect end_protected
