-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
XObI5BAuRGYhI+pqh//oJm46v/q9ALRHIOQVhZZM1XgFiMncrigGWt0PMm2iMry/72Aycz/RricR
MSK3DMxIBJWbhgMjR9PDN6VfqRW5ahm3Jwr/UNK3SIBBnX9RKkBeyGxpDFJjzDDFCQGe369LbLBh
ZrXMyRvOU4ARKcXEfj1mo0umjBIja4dNUUglWWzgelnYP7ZM0+ywVzV56IR32h12z4KTikPZptyY
qhtB2rdwf6xxtVZg/11+cq07n4Vm5pTNR8Qbnu61unG4j+WYY4uUNetwfmIsOOBXPthKtcOa8jYO
NeycCAaXo7rEi/jC0Ng5pUyD8xg9sbvvgxbHcQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5200)
`protect data_block
/44jNed06EXiLYdn7gELxDrPZcuVkmJNEsL3j04lNSEHOMYVP+ODR/ezbkonwBRJe0511gI/V4fw
O02qAgIiqjFSYtFxFSvdFnnegRh3mXKpX5xu9gnzoD7vDmpfCpuVso6ik0kgwXNqZX6OEZXCrolI
AoCSutmLWrXDDw7PHcdGS76kee83MePBGD7QKS2Z+rU+CHn+vULglVdW4oDVjZPA8NcpE9B9sOjX
kWeH4CjUxzZWGHY8PN1EouuyrhDRfgYEEev3ZdxP93fE+Q8ECJlvC3F4/ltGjJZtNy/jSkpk2DGe
BnQky7jF28dnFDvhkxwMWJOnUY+tjgqJsy1UB8vw52nrHUPkdhh5mxOOSHgsCmOXR9j6VmMK2Yg2
2XwR2jdXCiLqtnbMim7vfGbYgEe1Swq1WzQrzTVoOZF914W8qJ0MgDIjedOhsaF+pXpqmQ9Wpf2Z
z0g06DvoaciV2ONYhAN571aOOKQh/G0xfuzCQK8zHnugn8cpXxXu4pNlvQEcMVuyscAnOr8WtdsZ
HP4kDDUQBhyYwilByFavoFYKlKdHIQbHVl3CaODZli10BvEbUESOpI9b9Zik08KwppuwZnLV8FHP
oQgXNDonSpwtrGoiNS3uk4SRFMRTtXFYA6REd9PeZ7Tcmj5YoFLGdBJsZAwFYwX3XkS3RV4yYz3W
T74v7Hl68HZu45aYPPdAyQ8feECJ3gsoQLB7xoZvHRE1H9xF4ocLyCoWbcVNw6YgVPAvnQ/PcqHb
Qj4zfQkq0QZIKGAC2T1nu9UVg5ee8KMYyPhGfyOqZ67CVwCeskb2WsAij4RY0Ur/IVg0Ve8nuff9
O8AYyGvFRmTca8x9TAG97EhywsnkZPAHckRJSL0WPnZGPw5N87qnAcE/E5tolfblLTLZ37re7+hE
z4wXEekfhTFGl5jsWaU/nFJuVgi4v8Tj8RZI91GmvgzeEwjy30f0tSO0V2Mp/RO2Z+95TibSjNvs
hsnqacQWpNOgqJ/FP1tc257K+jo50m8e5nz0cV5t4zGk0NU3pfti3XATfDDtTgHrvn7JF34SNNMx
lSaAggIVpOvtOjmfx7NavocqZE6+ToAyWRUBVf28gygQ2qv2CyObe0Te5VgMkpAG8j5/dbyl0Eya
jQqF9QSyVS7U8PTMJwJJvyOsvRQY76Isy9p4sKc7WPK+LV3T6J2VERvz8QQsv7i+oF+P1ek+nU4y
DhePLARLMeCI3DJ48crIIseCXALvu1O7wAIqm+LKl8CnKafsG5c5WHIboh6IlEv2CU2HNndTpsxh
wKLZMSvQeXGO2fzUXlIozCb2BcxTmUjKevhUQJNCYjCjKlm6kE/WEiSR5kvb6oD8O4GOOsohRCuM
0tnpoPuooSF1XBjWbFs5fvyLJpo1R6y9SoeaxU8Horxb+VSjnJKBp21Zj8Ee+HwEDm60KgGtvrEz
XLYOOPGE/utFE9b8mvd2JKKp052jODuqDi6RczjszDwWcCN3lU0jteDv021Dp971lC6XyqQR7nq8
r5oxXlC7kEMkUijDmUFhAgNHov/HVXg4NAP91ftTOLuPdQ4mU+Y74jQW+po9DPbd39g0x1VlMHig
vO+iQ1wer3MoTd0zIGoy+6rVriu6pmOSrdVUGI8cDHvNV6CftR9m/dYKHB357SDp/Kap5dVIEhot
9T+QLePq0fsRGZOgHT5vaKwZySvWkrixMqhcaXcKqChhF+AITQ/3xoHsU0D7CWGt8g011M6kKeun
BhJQMtTnFZWxE/VXddS8pu1hUEj54aYA4AitSSZGGzZELvJyOugY3H62bu9eF0y47pOCL+IhnYDI
09pgDVre6h/81Ajgnii0Xtlugqml8nSXt8JxgfxB4tqYjla02EdILv9hTnWUNwQVO6uIGlgFkMXm
fbR1/6iFSub7fHM1I6YRLmwTNQUjHhDSO6bNsyBCzuv9/Ck4QKY+G3cHdkJenlepOmTKGaRlw8nM
K+QGZug4ZmAxUklFLJ/V0dVPd1vI7fmXEL7PkoiTCxupdwOmBjDI/0120IgVggr/TWO+Y2Iiv7Yx
Go/MlWReMoTAHXwkIjgcXSEcnxnhcRvAdw7DaX0nVihOvcymCY5fVSTUPnXJt5ghAF3NfdMgPeap
WYnYfL+5BK1p4vTAVCUGVLDtf16tMl72RAbVCtkq11sxrKbYHXVlWWr30kVdrJmlIL1l3g7bJDwx
RMrZeQfHMFESMXdQWgUrcpc1x0xBIu4FM9RdyZXBKCW+2FXUVEvI4p6XC1TCaLw5zkPL3pFX5eW6
MsdUdUqafh5mjoSZ8oYIXV2d+RamZ7n4HGJZ0lpiS6UFj0gAZADOdgmH+vz+TVokMqbHBJHjA4o/
wYTNogM/hMWJzML6u/IN/dM7ffuQkjGkN8JjKR33aHz0trNtYO7mOvOV3pZ4AYPR1xw12wTwuWYP
xbvO4MCNN8jro7Hzv8DzTP6UT86UTZDrCHPYvU+nUy2nO2oLUjCsfj/xfaWefTR1s12PLX2lBdp4
cleTMRIY4BjL7DCkxDYs/lioi/3Z/gTX0b08wg6rx3k7jtG1Cbt2uBggHb/DOIHQo8/p7S3Oi4do
Up9L+BcUsxm+VQsh80KykcLVXjuqESvvoCQX1WGJBO9ZI/I9V+zF4IimH2MAlBWNqZ+RYxj8n8ja
PYhiK+ggBw69jFROmazaUsySFIqU9aZrHXF67nt5s3jAGCJNgZcA58tnKFqKqoSsVbv5AaJqgwyp
AOTTwth/VprgfFhpCkAqVpvKwMB++iK2e71zLsREzlmIjXITvqnKd0FAf4/ZA9MABQElQKYoL1m2
tDEYqVCl/aqeZLsqK7eVY6e2z88YkwQLrdnQUJS7F9T60u4xZaf7PoaqrcZoTA16yT9L4JW+kAxN
Gj2PiDzuF+hzYs/xZroZlwDf1/FJnm0Tarvo1Ody9hNhg5rTlO4FyVHO0JRlyF2KcX/c29aIqTC4
Z482s9vHOJEeJCjBIeLYexvhgtoNGtdr7DmU1f3JytH7/ftYc5iUi0ZQ1t+0H5Bd0SNwQKsJwN4M
ICzx6hfF9/y/7+Xf68Cnyiw5+FO8gRgXQ2yzAJ2209DDU+EaQGIhwFI8xdqruWw/IJ8Qn02YXs3W
NM7lootLOZ6hrvvPko00UX1k14QHCyG0qnY+eK2b5VX9AkJbsxgdOrbxV4WsxEmUlmaUhZjETre3
19UldkCTG2Z8Stzb8FUdCLIQGB8V5E5oMntH/nc8urWm3dKvEgqZvNl/bLycV7Qr8BOVQLO+/XQ6
O0ydo1HuO2PHmDYMH8ooqIE8ZpL5sPqE6fSLcotrpaE1dJ6BRouQOdWJcJzBbvE/ItVouSlgJF2k
k04DtveRsuYkxRYje+jFQ821gbdBITJRVXx3/tk972Ksh/RD3OrOPTU72edMg/mWmHO92oRsVXic
576SPka45/eJtZmnzFW0s4lbuWB8rFHr9/TN8rH0M4wIghoJHPVX1z/lx10ovHgBPrn2DSRPqyPy
bqwpIvMGpqJztMuSDuCyRrncGbk97HYdpRpbwlfQSvVQlpt7AIccFjmU9gKzigYhEghL/l5bigwD
zP05gooOiTow6FJq6p7McAR1ENhdYVxlScyd3w9QTiHIdP4goT+onaNTEMOBjbqRNbfMOjcFZCvp
CzM52WexQa9Cl2VagHUkjAIP89BaAHtqMDQ8ea6DnzZjgPdfnIDtu9t1oFRXYtRBhvwGXGDzK8Rb
C/6n62ImDwpB76K5FjF/Fs1YU2RW9DOEk7O7g9y0iHUQ2u71ebiCz1MUoELrvKeusYcquqzQWbKk
32TbXaiJ7JQVfgD3yyKbcfRYO4qPpTJdflN6LZLG6Mq7eHJNvKVfly9uinvcKi1v18yxieXaoPPL
cOCN7qLbAZVeLcPmwehPa50zZdf6cK24LW3POTK+gGmPX+Mayc7FyLKE8qGxPcdbAt8bpdWTriUq
vg5Zb+UMtkPgluVQj3+pnGgyuJ7g/+j3eELxd3X3285K3bcm3FYGOda70Pf8cK+4SIcStfV4dctg
u3yw0VlKspG9UGyKmScn2WuG7rzaBugmMwk6mwGlJRT6LYtTw1u7oH3ljxzfek9iaNHfVH5zpRmu
HM/CF5njzIhs+tukPHgnFcpHDGL0O8k3CHrd3W0qS+LgXFEwHX6ShU1kdHsjgyIDpXW/eNOkzPcd
dUk8HD9DiPN2d6S6wY/r9WlK0Q36L5tHt8VYPJpUhNz5zZIJmIbDoZKL2YfxUwQ7DB9StdHnH7EU
c6KlwqRwzr/gJ05ZT2x0y3LqqoP+Iff7Ai9rIs3WELJCeBYvTX+dBz2sGtLfMDGlSrIPMouguND2
wElAWhVmkUeXvq22TBDD9CEDqGVPdXJ6QT2762PN9SrRFZi6QTmgJzJJxgXFbQa8Hd15x/zxZp1g
2Ry0L+sern/Bqu14e2pARSyiD0LAcS/5tXavoBjF4eJEJwXlNXauudSki7ninWrFHrJ46ByER3+J
cLA/c0/Sne0QhOQWwvMPkSxocBOF0SOI18PlcOcoFaNHoBv8OdfFR1rRg953gNe0N2AFXPQFQQbN
8HzwQH2X/dxsXU6FUB1puGCZAc+OotxQCcI1xlj/Om/wcdnghKfkZ4I/tB1hOOsm2RrJ52wYubnV
rv2k64slil/CMIEVM790iW8obg4mDz1E6wCHEHsWdybnIdvXtfYLgLx4aZqTO8cTwMCI+5nMyyFV
BWpPNxeOxyzjY5uHrGT058cEm+GW4ELO1luqgMF1NesZDKzowQxHkUKRW0n4ReXgQFjjgww+x5wW
W3b3v8oTJMViG2CvuNR16iwM16/W6ZWHTfL6kLTimBqPz0ixApfiCq4uvoxf6S5K3wdoC+o396HX
s3f0Pt6VYJfyX089BcOqHFS09zxVCuiRyDoSKmblkTN+dwGnahny+kyZTbIZokgQ+teTIPKpP/ff
IalmH0VMCbXEX/K2B++EsEqmdYI5QA6RB6s3OTTJBh8+4DwHpd3HNv3n+QRjb9B3i4GVZP72UB6C
mnMoKCvrepesGphcUGnboHLwYgehmPgBRr47rMlwMSIJkFL1JkhNY9488t5YqEs7C/1Tef1woRko
v2ujC2BZLdbxEjWvf+QU0Yyar6qt20Ewp5rF9TwJ47tbKQxcoPIjoT8bEITTJY5pKirQI8BVNiMd
NUBgNKZyrJtZjsy8aK/HKLC5EPJV9MrsrSN2nbgwgWgHLWArj+BG1ZLmT9pBjdV0x3mbS+lCQL9P
E/KYPA79Mmstwv2Wpyj+PYHKIlT1V0Tgbrc92KcRh3WpIOg32eoj6ND0r00Jjv8n/Oy/u6WboKDc
Uqhv3hpoo6tDti7lSaylhMfhqwlraPyJZSqkvp3gfqBfSq3hENQ2lYzMszd+/1L2TILPPuv8K69S
yeC1qCkOdVM92t4n7Kom01Rxd8wmCk9PqR6dc9TGIKtPfgnu9gTnTfYJHzo19ng62pxc9c3f+GyT
wxganndwQBg1HVBMREGqIPYbbdSH75aZmYzshBUYmrXJ17+Q4gqW2in8rPMtT/D0dfSTBMxmuXRK
fFXZyK/LGLZZHwxc9PmyXjZNcVCe3lWxhHHkMc+o9px1lYwfAR1N2+pHviNBbEj+uePADudM48yg
HWF+2AdJGR0+ADIzrBWN0ZJ1Dkeycx9g29z73es/GWgsT59A6Upn6yqM0855bVGWNWtbQsO7qQBC
sGx3EkBQSAZjrt62RM2JBtXhWau7knDuo+VNJ5lnSFQHW8xCQ1nAuaaWTDyFLtGJhghJgPJSigaK
PwYZFsNKUumAWg3daoG+TJ5fviY3EmFA7PVs8VtYtE8v08N19J1RZFSYkWTI9FFx1v7g4QbyKndT
w+KSqzrqM1OoRNXdaxdM9MjtZcka+VX1DL3E6j4TU6KqA3pfPbmdGJBCk3uqR7j0O/u3UJ0yVFvc
sN8mVBSzVAYlM1ZRamGu8e6RLBN8VGYDnfKD05Adzy8G89kMzPyyxJ3Bow9AIt7t2qm2tjnbM4cP
kJqjKdtPArmeutzKGQkYzpLnV3hvEoCMEF9oOIQiB3CGRnmU6nLF6AWFrZYuQkWF+QlAmyEVPuSg
w2+rU/oShu1Xk+o4v3rqNUY3RsE9HMdQwXHL8Q/GNxJ7K979eCx9YmF2JdvrFDoWyF56vi5mjqaR
alY0YFkWja8rpxuuNdP8vOgbTqtl+kGqx1JsOBys88wPTD0x9hPl3r5nLUfmmy3CcUVlswVw5jQH
Rdy9HiWSeUEqX/W278e+rriQ/W8ptOg+Aqv/1M/KHWRdqWZ+vF9Wyb7G0X9rfi8QfZumt+1ZEI3a
RAqc6lHICGU8mICiDutADKyxSAqbfYRko7ft8cR/x6bGVaEODyx9INLjcQW8nQ0/kvN0e+o9PU+j
lSSz/Zx6CtoHNGR1EznbVmDo8nJ1qG4gV2HsoblftmsDvznZqGDRGyqQRetgvBRvqKYYvj2yco/M
QDAbI3nlt7I7fJi5G+ygEJBwy5euqv+s95mPYp7LAbRNYD9BOAfdmDXiV9qC1nS7D2+lKfbGTAMg
HWIzcac7wzxPLXFk4XfN0LHLXhdpWI4k1us6B2eYnMAdOcbL3hteHyezXCWmQ0ze+LhylnJTmxry
NDgP6PXA7PLKsMi72F1FZtcc068Km/0FGGGN22WTt7pndAEyxMZ0Bng/UohkLLlc/qjjW2tW0AoU
didTwOXOclKARTjeETlh8m7SIqJUSX/Ki2ksUloSwwDSR9WHq80W3ikKE/4hpzqC5MQ0awRPcDaj
Kq4m5ockeohRXJST9gKQ1ycL/5720Pv2Alx3LfFzv1MlufGa1wNPx+8iZIs3yghu6+vPEI64SwaD
fA8TruwMKzYI/7gFx/cvDo9XVYYnrN8nYxwfYX50v8gfNMuz68QwNlnozJ+2tyvG3Bi2O3srpjyW
4/dNOjcAd0AZMP55fA==
`protect end_protected
