-- (C) 2001-2019 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 19.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
ahYvNnjoU8WFc/u2Yz522EFrQo/QG2qsZp1NQVnx3hF/kDwixdBojNOqSCgfyGP5
chES3uOp5mjsilaC6fWvocIp86i9ouxZJw5DMbYStjv4kPoyGr7UDvohQFd4r3yl
N5OBhU3+b6EZRiVMLte/At/w9ZlIotWGoNBrR0yRiak=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 2576)
`protect data_block
rNUeWlyraBsRSBh3021NPWZ9Wne0uTJP1qJNcHmtR7e2OjX6vxabPb4jVhJLWq6Q
jQRzEjp36nJ1Klm6cWoiJx3RTQSoxy5R4P/OkKej6g2sejCh2zpMRXHUrRJjcsNX
W7QECEEQPRTykNpxTlqhSB9rs035269p6VH5o1Bd+ZHOB7s7EekSno855nEN/zOZ
ddWyAv1NgnBLG1MgJaLdA/UGW1iNcpCKLdV+ROoiyl2pRNkvohmtci0vQnfYTMTM
jQ5KC3bA9gK+iT8ug4j0IeaBmtytx93QFNOXYmESms1CdJInTC+XNpBTACk1zjTt
r4pVgIB9eYwRo9YScEuVfN65zSwhqTPLLnvX2b1Oq63S2eUO/5nTdiZXqxx73dgI
WJ3GHBViia6RKMrQgaqQXRO05B2/HVSIbfxKACTdzCsneZ7+PzTzSCH9N+vwRWFU
02PYOVOtG4xq5rG3+2G9PTwSu09kN6FVsENEaqnz/LMHOn8jrAhNONCEnH4bMO9j
bXC8xMDSk8219096P5jyqCiQ22vyju5QPHfxSKi3u9Tug6XxbJoWneThwUSAdhTy
2ApPeIu550qBrJ+MTk8a77s+M5vmY2qLKRFp9b5EcQyBv8l3msWysbuKrdbCVOhn
Ysd7NKl2sfnwnuYxAJikOkXOYiOHmIsHsBasimnnhfIVzK21z/Wt7VU0FoUHWz7N
zqsXL7RHyP+4IBIimNNHkq7zuGEpYt+5Z6k9DYnT60ZhqjUFjsrBWrWC2RrzxEgI
j4HkyW0S8F7WQt0wtjpzIiRBhhFnBbWP90DMmMaxVGIt4AOmtHY5P84lVFNN973k
Vpm4jBs8KdF7BT8HByYZzWpF+5bSqO4LQY139CHRaMbhyOCVScHKiPovL0M8qt32
cxpe+2xlTNLNFtzdrxMKrqaV7ETXlPlEmPcK8KpbgonJCaZxrMlD2tOcsGcfA3bE
+c9vJrbHjpj+o1DVbUy8G+mRSMXQvb7gTjip8CM2GnRrTQ4dhue4H1VY1lnfA3JC
yHWrO7m5x+t5bqJEFd1F3CADsFJSiVpvTih0+Hc2m18dmRmewXQHfV0AaJqoKT6p
8I4kIYeO/gYOUIGV+MuxQF01lq21SWjyIt11renAGMn78n406iF1kqnNdVeyuRtl
TrXa4O/6+rz+NYrG2gFCPUF4yda3iqiMMR6sio+C5yEvzl2T10pow+T4mWTjWPZ6
lGZom1G49t0ovOkLu1uDrYCR/qohKhmf4giARVST/Q32DnH1GO3RBO/JTQKJJQ1P
m9Ds/xs43tkDYO+o55HuhoyURVAAPusvwGpX7FZRTxp21Bf61pf9B+KRqEkdvJ5r
WKJKfXu7eAds3UQUaTiehngGXWl2xs226cNv+wQ7cHiKGjjxg4pofwdgon2oUe4X
wyutZblZGRHvislqN3pyMn39eOcCWBqxxeIvri0puSrNf9vtODZQ0MAP7hVGULbm
tYQRdhIoDxOTMjpzXRJ95Yf0YN93o3EGxrB0lc8vQ5hjkSAx0W4FyFJ2KjHEJJ+p
tDni2VpYFmmaryfdEzpxp4uaXF5DemEwEEhHiJVCWOg/itnDqdD+YOOR+5DJeQJd
jjuV0ScVHja4u4jQlP0L38Ew8YCsTGzHkj/mek5UupMrMy6lKKtSmDOcrMroRSFb
J1Yz4MRNhXYmcNMlUq7g2SPj01t951D9MmcQDKtQODTBq03wbtAGzjOak7DF/jaz
PiPTgLEh/l5pCWOKhfbjOcYdFTPBzERrDeSSNxO0ixFDn9pvoyft4x4XTZfaLGsf
DRh2oY87V7Q5jXCgOovJZPnIf8JEv6UAAGikRDE0F0/pdc/l0FyNL9q1rW0Higlk
MJtx/KDSO5erpXUcYdQI5Dm1cgPffb+jXdnYk7qkCMAXYhSJU3QgKfB9fz2+ZYxK
+3vwnLUWx2FvlFPHEGD1WmwGmNxWtGyHilE2N2x1kgmc2D59S5AFkbbULxYGofYv
rJzIwgj2QH+TNzmLchktqpAt82vZ8WfGc+Ly0PEeTJc8MTQkbxqMjhThxYpMDSdm
PPcgra7nBPmJLHnxL2CkVgN4bMC0+37v4g6b5/cXI9WQuaMhBLteXUwb2ZjeycNh
7MkIbI67WV8ino2UeGpxD4pJtnz0DDEhyBQnER5WXWEo00iOWenWcrOll5Swk7CG
HnSRxw5rAhrwzEFfRsouSBLuAr4Ic+c9kEZ/rtxAcLamYKryf9hOJ9GuaasQ+DDv
6W2B4j4cRXboL2WjBzZ+ixIWzPM+1YNPPKi4J0wGjA99gfmoGUk2UM396tvQ7FJM
OI/tQX3Bkyv2Q+aZFa//cJrqMQJIxlZMHYpFlEDUHiZx05tcF+/c8E+taNxRs5VE
XSLy5BEbj7ezr3YNEtWD86xEY896n1WieBDxlLVyKaruFGGB94Sr43USjM4c1JFY
xHdpk0tJOa84hRzxmGlF9W7zGrf19NIpCN96YdqlWEJ07+/kQsuyYkzZMLMxcvTd
eQtOJeTcTbLRYvNWV9hht/2LDxc4xmb+biJiN9Yk3j4TJO66IRZNDEbYwBLZDlTy
r2pAe+U6QfqfGEB0IJl81iUc89r0p3muPKj6jZw0Uw2ImE8Ax8c4+BRH9BFS4qhm
ZyMNuysZ0/aVn5sGlDMEsvOO/9NU4YtlBhUU0uu1e3nmNk6KgQvA0CDgsZcelCZj
ndbr/UqKW5dEFhW2khZQKYE91GxMyXip9KfoXubpfyoXuaIsrcDqPiDUmeFHPYjY
q95DgmPTpG3ON1zib76hndeT5yBiCWrH/HwMjzE7O5JM7viY8O7RFBKKfIXxFDFz
LguHxQN5mFGlap+u3kaPpK1+kTJ5BtI5rJQAvZEB3tR4VpkhrHeWmnNFfy+qtUIR
ONwPe6vWsjR93AIUcuqXsH9W7n5SEHU9aVqdhfnfrMFTl54uw/jb+ec9n26KK1wE
kIPh0YVuMD+jFCqMNJBNc9qYBn9Vpk1KQqQ64m/M3FXuunemrCJioF1BuGld2raE
GLreQ0EzXCMRU3x3vmNd75+wcH8J7/fV3RQS/xc8QhxvESgb5lNaU2Z1ZZjJZRSr
Ohxusp7cEgrqVtyTqjGXca9qYYPXb2dCLpCXQhXNwNfe29zX/xY6Z9wTzu+FysXX
r9PwswnKnsEYytp5IEachSEf+xkylfYvXQY3PpqhPsEPZhDs+BiVg0h40/eEMpa0
1JdSQyorMeg2uzEfMCPDpk0YxlhBg1HQ2JP/aZSzQvRwbmaO36w/UhpM9zHfT9sV
1x2J1re9OZtdzplm/TUW+QMeW3frTzxJPrz9hW9oS7JTcKOnmK++hteCzFjXOkxJ
RmbcmZBMPWU9TLEGUeialnsTMiQuh4PFFdPHAX0/+H+Fhin1mVsoMUomTpsrGjD2
4tNo2mXespAjDg2ZCiOUKL0JXKGjaiptJ/FAWzHzr7o=
`protect end_protected
